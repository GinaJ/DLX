
module DLX ( Clk, Rst, exception );
  input Clk, Rst;
  output exception;
  wire   read_notWrite, \pipeline/Forward_sw1_mux ,
         \pipeline/regDst_to_mem[0] , \pipeline/regDst_to_mem[1] ,
         \pipeline/regDst_to_mem[3] , \pipeline/regDst_to_mem[4] ,
         \pipeline/MEM_controls_in_MEM[1] , \pipeline/WB_controls_in_MEMWB[0] ,
         \pipeline/WB_controls_in_MEMWB[1] ,
         \pipeline/MEM_controls_in_EXMEM[1] ,
         \pipeline/WB_controls_in_EXMEM[1] , \pipeline/WB_controls_in_IDEX[0] ,
         \pipeline/RegDst_to_WB[0] , \pipeline/RegDst_to_WB[1] ,
         \pipeline/RegDst_to_WB[2] , \pipeline/RegDst_to_WB[3] ,
         \pipeline/RegDst_to_WB[4] , \pipeline/EXE_controls_in_IDEX[0] ,
         \pipeline/EXE_controls_in_IDEX[1] ,
         \pipeline/EXE_controls_in_IDEX[2] ,
         \pipeline/EXE_controls_in_IDEX[3] ,
         \pipeline/EXE_controls_in_IDEX[4] ,
         \pipeline/EXE_controls_in_IDEX[5] ,
         \pipeline/EXE_controls_in_IDEX[6] ,
         \pipeline/EXE_controls_in_IDEX[7] ,
         \pipeline/EXE_controls_in_IDEX[8] , \pipeline/data_to_RF_from_WB[0] ,
         \pipeline/data_to_RF_from_WB[1] , \pipeline/data_to_RF_from_WB[2] ,
         \pipeline/data_to_RF_from_WB[3] , \pipeline/data_to_RF_from_WB[4] ,
         \pipeline/data_to_RF_from_WB[5] , \pipeline/data_to_RF_from_WB[6] ,
         \pipeline/data_to_RF_from_WB[7] , \pipeline/data_to_RF_from_WB[8] ,
         \pipeline/data_to_RF_from_WB[9] , \pipeline/data_to_RF_from_WB[10] ,
         \pipeline/data_to_RF_from_WB[11] , \pipeline/data_to_RF_from_WB[12] ,
         \pipeline/data_to_RF_from_WB[13] , \pipeline/data_to_RF_from_WB[14] ,
         \pipeline/data_to_RF_from_WB[15] , \pipeline/data_to_RF_from_WB[16] ,
         \pipeline/data_to_RF_from_WB[17] , \pipeline/data_to_RF_from_WB[18] ,
         \pipeline/data_to_RF_from_WB[19] , \pipeline/data_to_RF_from_WB[20] ,
         \pipeline/data_to_RF_from_WB[21] , \pipeline/data_to_RF_from_WB[22] ,
         \pipeline/data_to_RF_from_WB[23] , \pipeline/data_to_RF_from_WB[24] ,
         \pipeline/data_to_RF_from_WB[25] , \pipeline/data_to_RF_from_WB[26] ,
         \pipeline/data_to_RF_from_WB[27] , \pipeline/data_to_RF_from_WB[28] ,
         \pipeline/data_to_RF_from_WB[29] , \pipeline/data_to_RF_from_WB[30] ,
         \pipeline/data_to_RF_from_WB[31] , \pipeline/Alu_Out_Addr_to_mem[0] ,
         \pipeline/Alu_Out_Addr_to_mem[1] , \pipeline/Alu_Out_Addr_to_mem[2] ,
         \pipeline/Alu_Out_Addr_to_mem[3] , \pipeline/Alu_Out_Addr_to_mem[4] ,
         \pipeline/Alu_Out_Addr_to_mem[5] , \pipeline/Alu_Out_Addr_to_mem[6] ,
         \pipeline/Alu_Out_Addr_to_mem[7] , \pipeline/Alu_Out_Addr_to_mem[8] ,
         \pipeline/Alu_Out_Addr_to_mem[9] , \pipeline/Alu_Out_Addr_to_mem[10] ,
         \pipeline/Alu_Out_Addr_to_mem[11] ,
         \pipeline/Alu_Out_Addr_to_mem[12] ,
         \pipeline/Alu_Out_Addr_to_mem[13] ,
         \pipeline/Alu_Out_Addr_to_mem[14] ,
         \pipeline/Alu_Out_Addr_to_mem[15] ,
         \pipeline/Alu_Out_Addr_to_mem[16] ,
         \pipeline/Alu_Out_Addr_to_mem[17] ,
         \pipeline/Alu_Out_Addr_to_mem[18] ,
         \pipeline/Alu_Out_Addr_to_mem[19] ,
         \pipeline/Alu_Out_Addr_to_mem[20] ,
         \pipeline/Alu_Out_Addr_to_mem[21] ,
         \pipeline/Alu_Out_Addr_to_mem[22] ,
         \pipeline/Alu_Out_Addr_to_mem[23] ,
         \pipeline/Alu_Out_Addr_to_mem[24] ,
         \pipeline/Alu_Out_Addr_to_mem[25] ,
         \pipeline/Alu_Out_Addr_to_mem[26] ,
         \pipeline/Alu_Out_Addr_to_mem[27] ,
         \pipeline/Alu_Out_Addr_to_mem[28] ,
         \pipeline/Alu_Out_Addr_to_mem[29] ,
         \pipeline/Alu_Out_Addr_to_mem[30] ,
         \pipeline/Alu_Out_Addr_to_mem[31] , \pipeline/inst_IFID_DEC[26] ,
         \pipeline/inst_IFID_DEC[27] , \pipeline/inst_IFID_DEC[28] ,
         \pipeline/inst_IFID_DEC[29] , \pipeline/inst_IFID_DEC[30] ,
         \pipeline/inst_IFID_DEC[31] , \pipeline/nextPC_IFID_DEC[0] ,
         \pipeline/nextPC_IFID_DEC[1] , \pipeline/nextPC_IFID_DEC[2] ,
         \pipeline/nextPC_IFID_DEC[3] , \pipeline/nextPC_IFID_DEC[4] ,
         \pipeline/nextPC_IFID_DEC[5] , \pipeline/nextPC_IFID_DEC[6] ,
         \pipeline/nextPC_IFID_DEC[7] , \pipeline/nextPC_IFID_DEC[8] ,
         \pipeline/nextPC_IFID_DEC[9] , \pipeline/nextPC_IFID_DEC[10] ,
         \pipeline/nextPC_IFID_DEC[11] , \pipeline/nextPC_IFID_DEC[12] ,
         \pipeline/nextPC_IFID_DEC[13] , \pipeline/nextPC_IFID_DEC[14] ,
         \pipeline/nextPC_IFID_DEC[15] , \pipeline/nextPC_IFID_DEC[16] ,
         \pipeline/nextPC_IFID_DEC[17] , \pipeline/nextPC_IFID_DEC[18] ,
         \pipeline/nextPC_IFID_DEC[19] , \pipeline/nextPC_IFID_DEC[20] ,
         \pipeline/nextPC_IFID_DEC[21] , \pipeline/nextPC_IFID_DEC[22] ,
         \pipeline/nextPC_IFID_DEC[23] , \pipeline/nextPC_IFID_DEC[24] ,
         \pipeline/nextPC_IFID_DEC[25] , \pipeline/nextPC_IFID_DEC[26] ,
         \pipeline/nextPC_IFID_DEC[27] , \pipeline/nextPC_IFID_DEC[28] ,
         \pipeline/nextPC_IFID_DEC[29] , \pipeline/nextPC_IFID_DEC[30] ,
         \pipeline/stall , \pipeline/stageF/PC_plus4/N37 ,
         \pipeline/stageF/PC_plus4/N36 , \pipeline/stageF/PC_plus4/N35 ,
         \pipeline/stageF/PC_plus4/N34 , \pipeline/stageF/PC_plus4/N33 ,
         \pipeline/stageF/PC_plus4/N32 , \pipeline/stageF/PC_plus4/N31 ,
         \pipeline/stageF/PC_plus4/N30 , \pipeline/stageF/PC_plus4/N29 ,
         \pipeline/stageF/PC_plus4/N28 , \pipeline/stageF/PC_plus4/N27 ,
         \pipeline/stageF/PC_plus4/N26 , \pipeline/stageF/PC_plus4/N25 ,
         \pipeline/stageF/PC_plus4/N24 , \pipeline/stageF/PC_plus4/N23 ,
         \pipeline/stageF/PC_plus4/N22 , \pipeline/stageF/PC_plus4/N21 ,
         \pipeline/stageF/PC_plus4/N20 , \pipeline/stageF/PC_plus4/N19 ,
         \pipeline/stageF/PC_plus4/N18 , \pipeline/stageF/PC_plus4/N17 ,
         \pipeline/stageF/PC_plus4/N16 , \pipeline/stageF/PC_plus4/N15 ,
         \pipeline/stageF/PC_plus4/N14 , \pipeline/stageF/PC_plus4/N13 ,
         \pipeline/stageF/PC_plus4/N12 , \pipeline/stageF/PC_plus4/N11 ,
         \pipeline/stageF/PC_plus4/N10 , \pipeline/stageF/PC_plus4/N9 ,
         \pipeline/stageF/PC_reg/N31 , \pipeline/stageF/PC_reg/N30 ,
         \pipeline/stageF/PC_reg/N29 , \pipeline/stageF/PC_reg/N28 ,
         \pipeline/stageF/PC_reg/N27 , \pipeline/stageF/PC_reg/N26 ,
         \pipeline/stageF/PC_reg/N25 , \pipeline/stageF/PC_reg/N24 ,
         \pipeline/stageF/PC_reg/N23 , \pipeline/stageF/PC_reg/N22 ,
         \pipeline/stageF/PC_reg/N21 , \pipeline/stageF/PC_reg/N20 ,
         \pipeline/stageF/PC_reg/N19 , \pipeline/stageF/PC_reg/N18 ,
         \pipeline/stageF/PC_reg/N17 , \pipeline/stageF/PC_reg/N16 ,
         \pipeline/stageF/PC_reg/N15 , \pipeline/stageF/PC_reg/N14 ,
         \pipeline/stageF/PC_reg/N13 , \pipeline/stageF/PC_reg/N12 ,
         \pipeline/stageF/PC_reg/N11 , \pipeline/stageF/PC_reg/N10 ,
         \pipeline/stageF/PC_reg/N9 , \pipeline/stageF/PC_reg/N8 ,
         \pipeline/stageF/PC_reg/N7 , \pipeline/stageF/PC_reg/N6 ,
         \pipeline/stageF/PC_reg/N5 , \pipeline/stageF/PC_reg/N4 ,
         \pipeline/stageF/PC_reg/N3 , \pipeline/stageF/PC_reg/N2 ,
         \pipeline/stageF/PC_reg/N1 , \pipeline/stageF/PC_reg/N0 ,
         \pipeline/stageD/evaluate_jump_target/N63 ,
         \pipeline/stageD/evaluate_jump_target/N62 ,
         \pipeline/stageD/evaluate_jump_target/N61 ,
         \pipeline/stageD/evaluate_jump_target/N60 ,
         \pipeline/stageD/evaluate_jump_target/N59 ,
         \pipeline/stageD/evaluate_jump_target/N58 ,
         \pipeline/stageD/evaluate_jump_target/N57 ,
         \pipeline/stageD/evaluate_jump_target/N56 ,
         \pipeline/stageD/evaluate_jump_target/N55 ,
         \pipeline/stageD/evaluate_jump_target/N54 ,
         \pipeline/stageD/evaluate_jump_target/N53 ,
         \pipeline/stageD/evaluate_jump_target/N52 ,
         \pipeline/stageD/evaluate_jump_target/N51 ,
         \pipeline/stageD/evaluate_jump_target/N50 ,
         \pipeline/stageD/evaluate_jump_target/N49 ,
         \pipeline/stageD/evaluate_jump_target/N48 ,
         \pipeline/stageD/evaluate_jump_target/N47 ,
         \pipeline/stageD/evaluate_jump_target/N46 ,
         \pipeline/stageD/evaluate_jump_target/N45 ,
         \pipeline/stageD/evaluate_jump_target/N44 ,
         \pipeline/stageD/evaluate_jump_target/N43 ,
         \pipeline/stageD/evaluate_jump_target/N42 ,
         \pipeline/stageD/evaluate_jump_target/N41 ,
         \pipeline/stageD/evaluate_jump_target/N40 ,
         \pipeline/stageD/evaluate_jump_target/N39 ,
         \pipeline/stageD/evaluate_jump_target/N38 ,
         \pipeline/stageD/evaluate_jump_target/N37 ,
         \pipeline/stageD/evaluate_jump_target/N36 ,
         \pipeline/stageD/evaluate_jump_target/N35 ,
         \pipeline/stageD/evaluate_jump_target/N34 ,
         \pipeline/stageD/evaluate_jump_target/N33 ,
         \pipeline/RegFile_DEC_WB/RegBank[31][0] ,
         \pipeline/RegFile_DEC_WB/RegBank[31][1] ,
         \pipeline/RegFile_DEC_WB/RegBank[31][2] ,
         \pipeline/RegFile_DEC_WB/RegBank[31][3] ,
         \pipeline/RegFile_DEC_WB/RegBank[31][4] ,
         \pipeline/RegFile_DEC_WB/RegBank[31][5] ,
         \pipeline/RegFile_DEC_WB/RegBank[31][6] ,
         \pipeline/RegFile_DEC_WB/RegBank[31][7] ,
         \pipeline/RegFile_DEC_WB/RegBank[31][8] ,
         \pipeline/RegFile_DEC_WB/RegBank[31][9] ,
         \pipeline/RegFile_DEC_WB/RegBank[31][10] ,
         \pipeline/RegFile_DEC_WB/RegBank[31][11] ,
         \pipeline/RegFile_DEC_WB/RegBank[31][12] ,
         \pipeline/RegFile_DEC_WB/RegBank[31][13] ,
         \pipeline/RegFile_DEC_WB/RegBank[31][14] ,
         \pipeline/RegFile_DEC_WB/RegBank[31][15] ,
         \pipeline/RegFile_DEC_WB/RegBank[31][16] ,
         \pipeline/RegFile_DEC_WB/RegBank[31][17] ,
         \pipeline/RegFile_DEC_WB/RegBank[31][18] ,
         \pipeline/RegFile_DEC_WB/RegBank[31][19] ,
         \pipeline/RegFile_DEC_WB/RegBank[31][20] ,
         \pipeline/RegFile_DEC_WB/RegBank[31][21] ,
         \pipeline/RegFile_DEC_WB/RegBank[31][22] ,
         \pipeline/RegFile_DEC_WB/RegBank[31][23] ,
         \pipeline/RegFile_DEC_WB/RegBank[31][24] ,
         \pipeline/RegFile_DEC_WB/RegBank[31][25] ,
         \pipeline/RegFile_DEC_WB/RegBank[31][26] ,
         \pipeline/RegFile_DEC_WB/RegBank[31][27] ,
         \pipeline/RegFile_DEC_WB/RegBank[31][28] ,
         \pipeline/RegFile_DEC_WB/RegBank[31][29] ,
         \pipeline/RegFile_DEC_WB/RegBank[31][30] ,
         \pipeline/RegFile_DEC_WB/RegBank[31][31] ,
         \pipeline/RegFile_DEC_WB/RegBank[30][0] ,
         \pipeline/RegFile_DEC_WB/RegBank[30][1] ,
         \pipeline/RegFile_DEC_WB/RegBank[30][2] ,
         \pipeline/RegFile_DEC_WB/RegBank[30][3] ,
         \pipeline/RegFile_DEC_WB/RegBank[30][4] ,
         \pipeline/RegFile_DEC_WB/RegBank[30][5] ,
         \pipeline/RegFile_DEC_WB/RegBank[30][6] ,
         \pipeline/RegFile_DEC_WB/RegBank[30][7] ,
         \pipeline/RegFile_DEC_WB/RegBank[30][8] ,
         \pipeline/RegFile_DEC_WB/RegBank[30][9] ,
         \pipeline/RegFile_DEC_WB/RegBank[30][10] ,
         \pipeline/RegFile_DEC_WB/RegBank[30][11] ,
         \pipeline/RegFile_DEC_WB/RegBank[30][12] ,
         \pipeline/RegFile_DEC_WB/RegBank[30][13] ,
         \pipeline/RegFile_DEC_WB/RegBank[30][14] ,
         \pipeline/RegFile_DEC_WB/RegBank[30][15] ,
         \pipeline/RegFile_DEC_WB/RegBank[30][16] ,
         \pipeline/RegFile_DEC_WB/RegBank[30][17] ,
         \pipeline/RegFile_DEC_WB/RegBank[30][18] ,
         \pipeline/RegFile_DEC_WB/RegBank[30][19] ,
         \pipeline/RegFile_DEC_WB/RegBank[30][20] ,
         \pipeline/RegFile_DEC_WB/RegBank[30][21] ,
         \pipeline/RegFile_DEC_WB/RegBank[30][22] ,
         \pipeline/RegFile_DEC_WB/RegBank[30][23] ,
         \pipeline/RegFile_DEC_WB/RegBank[30][24] ,
         \pipeline/RegFile_DEC_WB/RegBank[30][25] ,
         \pipeline/RegFile_DEC_WB/RegBank[30][26] ,
         \pipeline/RegFile_DEC_WB/RegBank[30][27] ,
         \pipeline/RegFile_DEC_WB/RegBank[30][28] ,
         \pipeline/RegFile_DEC_WB/RegBank[30][29] ,
         \pipeline/RegFile_DEC_WB/RegBank[30][30] ,
         \pipeline/RegFile_DEC_WB/RegBank[30][31] ,
         \pipeline/RegFile_DEC_WB/RegBank[29][0] ,
         \pipeline/RegFile_DEC_WB/RegBank[29][1] ,
         \pipeline/RegFile_DEC_WB/RegBank[29][2] ,
         \pipeline/RegFile_DEC_WB/RegBank[29][3] ,
         \pipeline/RegFile_DEC_WB/RegBank[29][4] ,
         \pipeline/RegFile_DEC_WB/RegBank[29][5] ,
         \pipeline/RegFile_DEC_WB/RegBank[29][6] ,
         \pipeline/RegFile_DEC_WB/RegBank[29][7] ,
         \pipeline/RegFile_DEC_WB/RegBank[29][8] ,
         \pipeline/RegFile_DEC_WB/RegBank[29][9] ,
         \pipeline/RegFile_DEC_WB/RegBank[29][10] ,
         \pipeline/RegFile_DEC_WB/RegBank[29][11] ,
         \pipeline/RegFile_DEC_WB/RegBank[29][12] ,
         \pipeline/RegFile_DEC_WB/RegBank[29][13] ,
         \pipeline/RegFile_DEC_WB/RegBank[29][14] ,
         \pipeline/RegFile_DEC_WB/RegBank[29][15] ,
         \pipeline/RegFile_DEC_WB/RegBank[29][16] ,
         \pipeline/RegFile_DEC_WB/RegBank[29][17] ,
         \pipeline/RegFile_DEC_WB/RegBank[29][18] ,
         \pipeline/RegFile_DEC_WB/RegBank[29][19] ,
         \pipeline/RegFile_DEC_WB/RegBank[29][20] ,
         \pipeline/RegFile_DEC_WB/RegBank[29][21] ,
         \pipeline/RegFile_DEC_WB/RegBank[29][22] ,
         \pipeline/RegFile_DEC_WB/RegBank[29][23] ,
         \pipeline/RegFile_DEC_WB/RegBank[29][24] ,
         \pipeline/RegFile_DEC_WB/RegBank[29][25] ,
         \pipeline/RegFile_DEC_WB/RegBank[29][26] ,
         \pipeline/RegFile_DEC_WB/RegBank[29][27] ,
         \pipeline/RegFile_DEC_WB/RegBank[29][28] ,
         \pipeline/RegFile_DEC_WB/RegBank[29][29] ,
         \pipeline/RegFile_DEC_WB/RegBank[29][30] ,
         \pipeline/RegFile_DEC_WB/RegBank[29][31] ,
         \pipeline/RegFile_DEC_WB/RegBank[28][0] ,
         \pipeline/RegFile_DEC_WB/RegBank[28][1] ,
         \pipeline/RegFile_DEC_WB/RegBank[28][2] ,
         \pipeline/RegFile_DEC_WB/RegBank[28][3] ,
         \pipeline/RegFile_DEC_WB/RegBank[28][4] ,
         \pipeline/RegFile_DEC_WB/RegBank[28][5] ,
         \pipeline/RegFile_DEC_WB/RegBank[28][6] ,
         \pipeline/RegFile_DEC_WB/RegBank[28][7] ,
         \pipeline/RegFile_DEC_WB/RegBank[28][8] ,
         \pipeline/RegFile_DEC_WB/RegBank[28][9] ,
         \pipeline/RegFile_DEC_WB/RegBank[28][10] ,
         \pipeline/RegFile_DEC_WB/RegBank[28][11] ,
         \pipeline/RegFile_DEC_WB/RegBank[28][12] ,
         \pipeline/RegFile_DEC_WB/RegBank[28][13] ,
         \pipeline/RegFile_DEC_WB/RegBank[28][14] ,
         \pipeline/RegFile_DEC_WB/RegBank[28][15] ,
         \pipeline/RegFile_DEC_WB/RegBank[28][16] ,
         \pipeline/RegFile_DEC_WB/RegBank[28][17] ,
         \pipeline/RegFile_DEC_WB/RegBank[28][18] ,
         \pipeline/RegFile_DEC_WB/RegBank[28][19] ,
         \pipeline/RegFile_DEC_WB/RegBank[28][20] ,
         \pipeline/RegFile_DEC_WB/RegBank[28][21] ,
         \pipeline/RegFile_DEC_WB/RegBank[28][22] ,
         \pipeline/RegFile_DEC_WB/RegBank[28][23] ,
         \pipeline/RegFile_DEC_WB/RegBank[28][24] ,
         \pipeline/RegFile_DEC_WB/RegBank[28][25] ,
         \pipeline/RegFile_DEC_WB/RegBank[28][26] ,
         \pipeline/RegFile_DEC_WB/RegBank[28][27] ,
         \pipeline/RegFile_DEC_WB/RegBank[28][28] ,
         \pipeline/RegFile_DEC_WB/RegBank[28][29] ,
         \pipeline/RegFile_DEC_WB/RegBank[28][30] ,
         \pipeline/RegFile_DEC_WB/RegBank[28][31] ,
         \pipeline/RegFile_DEC_WB/RegBank[27][0] ,
         \pipeline/RegFile_DEC_WB/RegBank[27][1] ,
         \pipeline/RegFile_DEC_WB/RegBank[27][2] ,
         \pipeline/RegFile_DEC_WB/RegBank[27][3] ,
         \pipeline/RegFile_DEC_WB/RegBank[27][4] ,
         \pipeline/RegFile_DEC_WB/RegBank[27][5] ,
         \pipeline/RegFile_DEC_WB/RegBank[27][6] ,
         \pipeline/RegFile_DEC_WB/RegBank[27][7] ,
         \pipeline/RegFile_DEC_WB/RegBank[27][8] ,
         \pipeline/RegFile_DEC_WB/RegBank[27][9] ,
         \pipeline/RegFile_DEC_WB/RegBank[27][10] ,
         \pipeline/RegFile_DEC_WB/RegBank[27][11] ,
         \pipeline/RegFile_DEC_WB/RegBank[27][12] ,
         \pipeline/RegFile_DEC_WB/RegBank[27][13] ,
         \pipeline/RegFile_DEC_WB/RegBank[27][14] ,
         \pipeline/RegFile_DEC_WB/RegBank[27][15] ,
         \pipeline/RegFile_DEC_WB/RegBank[27][16] ,
         \pipeline/RegFile_DEC_WB/RegBank[27][17] ,
         \pipeline/RegFile_DEC_WB/RegBank[27][18] ,
         \pipeline/RegFile_DEC_WB/RegBank[27][19] ,
         \pipeline/RegFile_DEC_WB/RegBank[27][20] ,
         \pipeline/RegFile_DEC_WB/RegBank[27][21] ,
         \pipeline/RegFile_DEC_WB/RegBank[27][22] ,
         \pipeline/RegFile_DEC_WB/RegBank[27][23] ,
         \pipeline/RegFile_DEC_WB/RegBank[27][24] ,
         \pipeline/RegFile_DEC_WB/RegBank[27][25] ,
         \pipeline/RegFile_DEC_WB/RegBank[27][26] ,
         \pipeline/RegFile_DEC_WB/RegBank[27][27] ,
         \pipeline/RegFile_DEC_WB/RegBank[27][28] ,
         \pipeline/RegFile_DEC_WB/RegBank[27][29] ,
         \pipeline/RegFile_DEC_WB/RegBank[27][30] ,
         \pipeline/RegFile_DEC_WB/RegBank[27][31] ,
         \pipeline/RegFile_DEC_WB/RegBank[26][0] ,
         \pipeline/RegFile_DEC_WB/RegBank[26][1] ,
         \pipeline/RegFile_DEC_WB/RegBank[26][2] ,
         \pipeline/RegFile_DEC_WB/RegBank[26][3] ,
         \pipeline/RegFile_DEC_WB/RegBank[26][4] ,
         \pipeline/RegFile_DEC_WB/RegBank[26][5] ,
         \pipeline/RegFile_DEC_WB/RegBank[26][6] ,
         \pipeline/RegFile_DEC_WB/RegBank[26][7] ,
         \pipeline/RegFile_DEC_WB/RegBank[26][8] ,
         \pipeline/RegFile_DEC_WB/RegBank[26][9] ,
         \pipeline/RegFile_DEC_WB/RegBank[26][10] ,
         \pipeline/RegFile_DEC_WB/RegBank[26][11] ,
         \pipeline/RegFile_DEC_WB/RegBank[26][12] ,
         \pipeline/RegFile_DEC_WB/RegBank[26][13] ,
         \pipeline/RegFile_DEC_WB/RegBank[26][14] ,
         \pipeline/RegFile_DEC_WB/RegBank[26][15] ,
         \pipeline/RegFile_DEC_WB/RegBank[26][16] ,
         \pipeline/RegFile_DEC_WB/RegBank[26][17] ,
         \pipeline/RegFile_DEC_WB/RegBank[26][18] ,
         \pipeline/RegFile_DEC_WB/RegBank[26][19] ,
         \pipeline/RegFile_DEC_WB/RegBank[26][20] ,
         \pipeline/RegFile_DEC_WB/RegBank[26][21] ,
         \pipeline/RegFile_DEC_WB/RegBank[26][22] ,
         \pipeline/RegFile_DEC_WB/RegBank[26][23] ,
         \pipeline/RegFile_DEC_WB/RegBank[26][24] ,
         \pipeline/RegFile_DEC_WB/RegBank[26][25] ,
         \pipeline/RegFile_DEC_WB/RegBank[26][26] ,
         \pipeline/RegFile_DEC_WB/RegBank[26][27] ,
         \pipeline/RegFile_DEC_WB/RegBank[26][28] ,
         \pipeline/RegFile_DEC_WB/RegBank[26][29] ,
         \pipeline/RegFile_DEC_WB/RegBank[26][30] ,
         \pipeline/RegFile_DEC_WB/RegBank[26][31] ,
         \pipeline/RegFile_DEC_WB/RegBank[25][0] ,
         \pipeline/RegFile_DEC_WB/RegBank[25][1] ,
         \pipeline/RegFile_DEC_WB/RegBank[25][2] ,
         \pipeline/RegFile_DEC_WB/RegBank[25][3] ,
         \pipeline/RegFile_DEC_WB/RegBank[25][4] ,
         \pipeline/RegFile_DEC_WB/RegBank[25][5] ,
         \pipeline/RegFile_DEC_WB/RegBank[25][6] ,
         \pipeline/RegFile_DEC_WB/RegBank[25][7] ,
         \pipeline/RegFile_DEC_WB/RegBank[25][8] ,
         \pipeline/RegFile_DEC_WB/RegBank[25][9] ,
         \pipeline/RegFile_DEC_WB/RegBank[25][10] ,
         \pipeline/RegFile_DEC_WB/RegBank[25][11] ,
         \pipeline/RegFile_DEC_WB/RegBank[25][12] ,
         \pipeline/RegFile_DEC_WB/RegBank[25][13] ,
         \pipeline/RegFile_DEC_WB/RegBank[25][14] ,
         \pipeline/RegFile_DEC_WB/RegBank[25][15] ,
         \pipeline/RegFile_DEC_WB/RegBank[25][16] ,
         \pipeline/RegFile_DEC_WB/RegBank[25][17] ,
         \pipeline/RegFile_DEC_WB/RegBank[25][18] ,
         \pipeline/RegFile_DEC_WB/RegBank[25][19] ,
         \pipeline/RegFile_DEC_WB/RegBank[25][20] ,
         \pipeline/RegFile_DEC_WB/RegBank[25][21] ,
         \pipeline/RegFile_DEC_WB/RegBank[25][22] ,
         \pipeline/RegFile_DEC_WB/RegBank[25][23] ,
         \pipeline/RegFile_DEC_WB/RegBank[25][24] ,
         \pipeline/RegFile_DEC_WB/RegBank[25][25] ,
         \pipeline/RegFile_DEC_WB/RegBank[25][26] ,
         \pipeline/RegFile_DEC_WB/RegBank[25][27] ,
         \pipeline/RegFile_DEC_WB/RegBank[25][28] ,
         \pipeline/RegFile_DEC_WB/RegBank[25][29] ,
         \pipeline/RegFile_DEC_WB/RegBank[25][30] ,
         \pipeline/RegFile_DEC_WB/RegBank[25][31] ,
         \pipeline/RegFile_DEC_WB/RegBank[24][0] ,
         \pipeline/RegFile_DEC_WB/RegBank[24][1] ,
         \pipeline/RegFile_DEC_WB/RegBank[24][2] ,
         \pipeline/RegFile_DEC_WB/RegBank[24][3] ,
         \pipeline/RegFile_DEC_WB/RegBank[24][4] ,
         \pipeline/RegFile_DEC_WB/RegBank[24][5] ,
         \pipeline/RegFile_DEC_WB/RegBank[24][6] ,
         \pipeline/RegFile_DEC_WB/RegBank[24][7] ,
         \pipeline/RegFile_DEC_WB/RegBank[24][8] ,
         \pipeline/RegFile_DEC_WB/RegBank[24][9] ,
         \pipeline/RegFile_DEC_WB/RegBank[24][10] ,
         \pipeline/RegFile_DEC_WB/RegBank[24][11] ,
         \pipeline/RegFile_DEC_WB/RegBank[24][12] ,
         \pipeline/RegFile_DEC_WB/RegBank[24][13] ,
         \pipeline/RegFile_DEC_WB/RegBank[24][14] ,
         \pipeline/RegFile_DEC_WB/RegBank[24][15] ,
         \pipeline/RegFile_DEC_WB/RegBank[24][16] ,
         \pipeline/RegFile_DEC_WB/RegBank[24][17] ,
         \pipeline/RegFile_DEC_WB/RegBank[24][18] ,
         \pipeline/RegFile_DEC_WB/RegBank[24][19] ,
         \pipeline/RegFile_DEC_WB/RegBank[24][20] ,
         \pipeline/RegFile_DEC_WB/RegBank[24][21] ,
         \pipeline/RegFile_DEC_WB/RegBank[24][22] ,
         \pipeline/RegFile_DEC_WB/RegBank[24][23] ,
         \pipeline/RegFile_DEC_WB/RegBank[24][24] ,
         \pipeline/RegFile_DEC_WB/RegBank[24][25] ,
         \pipeline/RegFile_DEC_WB/RegBank[24][26] ,
         \pipeline/RegFile_DEC_WB/RegBank[24][27] ,
         \pipeline/RegFile_DEC_WB/RegBank[24][28] ,
         \pipeline/RegFile_DEC_WB/RegBank[24][29] ,
         \pipeline/RegFile_DEC_WB/RegBank[24][30] ,
         \pipeline/RegFile_DEC_WB/RegBank[24][31] ,
         \pipeline/RegFile_DEC_WB/RegBank[23][0] ,
         \pipeline/RegFile_DEC_WB/RegBank[23][1] ,
         \pipeline/RegFile_DEC_WB/RegBank[23][2] ,
         \pipeline/RegFile_DEC_WB/RegBank[23][3] ,
         \pipeline/RegFile_DEC_WB/RegBank[23][4] ,
         \pipeline/RegFile_DEC_WB/RegBank[23][5] ,
         \pipeline/RegFile_DEC_WB/RegBank[23][6] ,
         \pipeline/RegFile_DEC_WB/RegBank[23][7] ,
         \pipeline/RegFile_DEC_WB/RegBank[23][8] ,
         \pipeline/RegFile_DEC_WB/RegBank[23][9] ,
         \pipeline/RegFile_DEC_WB/RegBank[23][10] ,
         \pipeline/RegFile_DEC_WB/RegBank[23][11] ,
         \pipeline/RegFile_DEC_WB/RegBank[23][12] ,
         \pipeline/RegFile_DEC_WB/RegBank[23][13] ,
         \pipeline/RegFile_DEC_WB/RegBank[23][14] ,
         \pipeline/RegFile_DEC_WB/RegBank[23][15] ,
         \pipeline/RegFile_DEC_WB/RegBank[23][16] ,
         \pipeline/RegFile_DEC_WB/RegBank[23][17] ,
         \pipeline/RegFile_DEC_WB/RegBank[23][18] ,
         \pipeline/RegFile_DEC_WB/RegBank[23][19] ,
         \pipeline/RegFile_DEC_WB/RegBank[23][20] ,
         \pipeline/RegFile_DEC_WB/RegBank[23][21] ,
         \pipeline/RegFile_DEC_WB/RegBank[23][22] ,
         \pipeline/RegFile_DEC_WB/RegBank[23][23] ,
         \pipeline/RegFile_DEC_WB/RegBank[23][24] ,
         \pipeline/RegFile_DEC_WB/RegBank[23][25] ,
         \pipeline/RegFile_DEC_WB/RegBank[23][26] ,
         \pipeline/RegFile_DEC_WB/RegBank[23][27] ,
         \pipeline/RegFile_DEC_WB/RegBank[23][28] ,
         \pipeline/RegFile_DEC_WB/RegBank[23][29] ,
         \pipeline/RegFile_DEC_WB/RegBank[23][30] ,
         \pipeline/RegFile_DEC_WB/RegBank[23][31] ,
         \pipeline/RegFile_DEC_WB/RegBank[22][0] ,
         \pipeline/RegFile_DEC_WB/RegBank[22][1] ,
         \pipeline/RegFile_DEC_WB/RegBank[22][2] ,
         \pipeline/RegFile_DEC_WB/RegBank[22][3] ,
         \pipeline/RegFile_DEC_WB/RegBank[22][4] ,
         \pipeline/RegFile_DEC_WB/RegBank[22][5] ,
         \pipeline/RegFile_DEC_WB/RegBank[22][6] ,
         \pipeline/RegFile_DEC_WB/RegBank[22][7] ,
         \pipeline/RegFile_DEC_WB/RegBank[22][8] ,
         \pipeline/RegFile_DEC_WB/RegBank[22][9] ,
         \pipeline/RegFile_DEC_WB/RegBank[22][10] ,
         \pipeline/RegFile_DEC_WB/RegBank[22][11] ,
         \pipeline/RegFile_DEC_WB/RegBank[22][12] ,
         \pipeline/RegFile_DEC_WB/RegBank[22][13] ,
         \pipeline/RegFile_DEC_WB/RegBank[22][14] ,
         \pipeline/RegFile_DEC_WB/RegBank[22][15] ,
         \pipeline/RegFile_DEC_WB/RegBank[22][16] ,
         \pipeline/RegFile_DEC_WB/RegBank[22][17] ,
         \pipeline/RegFile_DEC_WB/RegBank[22][18] ,
         \pipeline/RegFile_DEC_WB/RegBank[22][19] ,
         \pipeline/RegFile_DEC_WB/RegBank[22][20] ,
         \pipeline/RegFile_DEC_WB/RegBank[22][21] ,
         \pipeline/RegFile_DEC_WB/RegBank[22][22] ,
         \pipeline/RegFile_DEC_WB/RegBank[22][23] ,
         \pipeline/RegFile_DEC_WB/RegBank[22][24] ,
         \pipeline/RegFile_DEC_WB/RegBank[22][25] ,
         \pipeline/RegFile_DEC_WB/RegBank[22][26] ,
         \pipeline/RegFile_DEC_WB/RegBank[22][27] ,
         \pipeline/RegFile_DEC_WB/RegBank[22][28] ,
         \pipeline/RegFile_DEC_WB/RegBank[22][29] ,
         \pipeline/RegFile_DEC_WB/RegBank[22][30] ,
         \pipeline/RegFile_DEC_WB/RegBank[22][31] ,
         \pipeline/RegFile_DEC_WB/RegBank[21][0] ,
         \pipeline/RegFile_DEC_WB/RegBank[21][1] ,
         \pipeline/RegFile_DEC_WB/RegBank[21][2] ,
         \pipeline/RegFile_DEC_WB/RegBank[21][3] ,
         \pipeline/RegFile_DEC_WB/RegBank[21][4] ,
         \pipeline/RegFile_DEC_WB/RegBank[21][5] ,
         \pipeline/RegFile_DEC_WB/RegBank[21][6] ,
         \pipeline/RegFile_DEC_WB/RegBank[21][7] ,
         \pipeline/RegFile_DEC_WB/RegBank[21][8] ,
         \pipeline/RegFile_DEC_WB/RegBank[21][9] ,
         \pipeline/RegFile_DEC_WB/RegBank[21][10] ,
         \pipeline/RegFile_DEC_WB/RegBank[21][11] ,
         \pipeline/RegFile_DEC_WB/RegBank[21][12] ,
         \pipeline/RegFile_DEC_WB/RegBank[21][13] ,
         \pipeline/RegFile_DEC_WB/RegBank[21][14] ,
         \pipeline/RegFile_DEC_WB/RegBank[21][15] ,
         \pipeline/RegFile_DEC_WB/RegBank[21][16] ,
         \pipeline/RegFile_DEC_WB/RegBank[21][17] ,
         \pipeline/RegFile_DEC_WB/RegBank[21][18] ,
         \pipeline/RegFile_DEC_WB/RegBank[21][19] ,
         \pipeline/RegFile_DEC_WB/RegBank[21][20] ,
         \pipeline/RegFile_DEC_WB/RegBank[21][21] ,
         \pipeline/RegFile_DEC_WB/RegBank[21][22] ,
         \pipeline/RegFile_DEC_WB/RegBank[21][23] ,
         \pipeline/RegFile_DEC_WB/RegBank[21][24] ,
         \pipeline/RegFile_DEC_WB/RegBank[21][25] ,
         \pipeline/RegFile_DEC_WB/RegBank[21][26] ,
         \pipeline/RegFile_DEC_WB/RegBank[21][27] ,
         \pipeline/RegFile_DEC_WB/RegBank[21][28] ,
         \pipeline/RegFile_DEC_WB/RegBank[21][29] ,
         \pipeline/RegFile_DEC_WB/RegBank[21][30] ,
         \pipeline/RegFile_DEC_WB/RegBank[21][31] ,
         \pipeline/RegFile_DEC_WB/RegBank[20][0] ,
         \pipeline/RegFile_DEC_WB/RegBank[20][1] ,
         \pipeline/RegFile_DEC_WB/RegBank[20][2] ,
         \pipeline/RegFile_DEC_WB/RegBank[20][3] ,
         \pipeline/RegFile_DEC_WB/RegBank[20][4] ,
         \pipeline/RegFile_DEC_WB/RegBank[20][5] ,
         \pipeline/RegFile_DEC_WB/RegBank[20][6] ,
         \pipeline/RegFile_DEC_WB/RegBank[20][7] ,
         \pipeline/RegFile_DEC_WB/RegBank[20][8] ,
         \pipeline/RegFile_DEC_WB/RegBank[20][9] ,
         \pipeline/RegFile_DEC_WB/RegBank[20][10] ,
         \pipeline/RegFile_DEC_WB/RegBank[20][11] ,
         \pipeline/RegFile_DEC_WB/RegBank[20][12] ,
         \pipeline/RegFile_DEC_WB/RegBank[20][13] ,
         \pipeline/RegFile_DEC_WB/RegBank[20][14] ,
         \pipeline/RegFile_DEC_WB/RegBank[20][15] ,
         \pipeline/RegFile_DEC_WB/RegBank[20][16] ,
         \pipeline/RegFile_DEC_WB/RegBank[20][17] ,
         \pipeline/RegFile_DEC_WB/RegBank[20][18] ,
         \pipeline/RegFile_DEC_WB/RegBank[20][19] ,
         \pipeline/RegFile_DEC_WB/RegBank[20][20] ,
         \pipeline/RegFile_DEC_WB/RegBank[20][21] ,
         \pipeline/RegFile_DEC_WB/RegBank[20][22] ,
         \pipeline/RegFile_DEC_WB/RegBank[20][23] ,
         \pipeline/RegFile_DEC_WB/RegBank[20][24] ,
         \pipeline/RegFile_DEC_WB/RegBank[20][25] ,
         \pipeline/RegFile_DEC_WB/RegBank[20][26] ,
         \pipeline/RegFile_DEC_WB/RegBank[20][27] ,
         \pipeline/RegFile_DEC_WB/RegBank[20][28] ,
         \pipeline/RegFile_DEC_WB/RegBank[20][29] ,
         \pipeline/RegFile_DEC_WB/RegBank[20][30] ,
         \pipeline/RegFile_DEC_WB/RegBank[20][31] ,
         \pipeline/RegFile_DEC_WB/RegBank[19][0] ,
         \pipeline/RegFile_DEC_WB/RegBank[19][1] ,
         \pipeline/RegFile_DEC_WB/RegBank[19][2] ,
         \pipeline/RegFile_DEC_WB/RegBank[19][3] ,
         \pipeline/RegFile_DEC_WB/RegBank[19][4] ,
         \pipeline/RegFile_DEC_WB/RegBank[19][5] ,
         \pipeline/RegFile_DEC_WB/RegBank[19][6] ,
         \pipeline/RegFile_DEC_WB/RegBank[19][7] ,
         \pipeline/RegFile_DEC_WB/RegBank[19][8] ,
         \pipeline/RegFile_DEC_WB/RegBank[19][9] ,
         \pipeline/RegFile_DEC_WB/RegBank[19][10] ,
         \pipeline/RegFile_DEC_WB/RegBank[19][11] ,
         \pipeline/RegFile_DEC_WB/RegBank[19][12] ,
         \pipeline/RegFile_DEC_WB/RegBank[19][13] ,
         \pipeline/RegFile_DEC_WB/RegBank[19][14] ,
         \pipeline/RegFile_DEC_WB/RegBank[19][15] ,
         \pipeline/RegFile_DEC_WB/RegBank[19][16] ,
         \pipeline/RegFile_DEC_WB/RegBank[19][17] ,
         \pipeline/RegFile_DEC_WB/RegBank[19][18] ,
         \pipeline/RegFile_DEC_WB/RegBank[19][19] ,
         \pipeline/RegFile_DEC_WB/RegBank[19][20] ,
         \pipeline/RegFile_DEC_WB/RegBank[19][21] ,
         \pipeline/RegFile_DEC_WB/RegBank[19][22] ,
         \pipeline/RegFile_DEC_WB/RegBank[19][23] ,
         \pipeline/RegFile_DEC_WB/RegBank[19][24] ,
         \pipeline/RegFile_DEC_WB/RegBank[19][25] ,
         \pipeline/RegFile_DEC_WB/RegBank[19][26] ,
         \pipeline/RegFile_DEC_WB/RegBank[19][27] ,
         \pipeline/RegFile_DEC_WB/RegBank[19][28] ,
         \pipeline/RegFile_DEC_WB/RegBank[19][29] ,
         \pipeline/RegFile_DEC_WB/RegBank[19][30] ,
         \pipeline/RegFile_DEC_WB/RegBank[19][31] ,
         \pipeline/RegFile_DEC_WB/RegBank[18][0] ,
         \pipeline/RegFile_DEC_WB/RegBank[18][1] ,
         \pipeline/RegFile_DEC_WB/RegBank[18][2] ,
         \pipeline/RegFile_DEC_WB/RegBank[18][3] ,
         \pipeline/RegFile_DEC_WB/RegBank[18][4] ,
         \pipeline/RegFile_DEC_WB/RegBank[18][5] ,
         \pipeline/RegFile_DEC_WB/RegBank[18][6] ,
         \pipeline/RegFile_DEC_WB/RegBank[18][7] ,
         \pipeline/RegFile_DEC_WB/RegBank[18][8] ,
         \pipeline/RegFile_DEC_WB/RegBank[18][9] ,
         \pipeline/RegFile_DEC_WB/RegBank[18][10] ,
         \pipeline/RegFile_DEC_WB/RegBank[18][11] ,
         \pipeline/RegFile_DEC_WB/RegBank[18][12] ,
         \pipeline/RegFile_DEC_WB/RegBank[18][13] ,
         \pipeline/RegFile_DEC_WB/RegBank[18][14] ,
         \pipeline/RegFile_DEC_WB/RegBank[18][15] ,
         \pipeline/RegFile_DEC_WB/RegBank[18][16] ,
         \pipeline/RegFile_DEC_WB/RegBank[18][17] ,
         \pipeline/RegFile_DEC_WB/RegBank[18][18] ,
         \pipeline/RegFile_DEC_WB/RegBank[18][19] ,
         \pipeline/RegFile_DEC_WB/RegBank[18][20] ,
         \pipeline/RegFile_DEC_WB/RegBank[18][21] ,
         \pipeline/RegFile_DEC_WB/RegBank[18][22] ,
         \pipeline/RegFile_DEC_WB/RegBank[18][23] ,
         \pipeline/RegFile_DEC_WB/RegBank[18][24] ,
         \pipeline/RegFile_DEC_WB/RegBank[18][25] ,
         \pipeline/RegFile_DEC_WB/RegBank[18][26] ,
         \pipeline/RegFile_DEC_WB/RegBank[18][27] ,
         \pipeline/RegFile_DEC_WB/RegBank[18][28] ,
         \pipeline/RegFile_DEC_WB/RegBank[18][29] ,
         \pipeline/RegFile_DEC_WB/RegBank[18][30] ,
         \pipeline/RegFile_DEC_WB/RegBank[18][31] ,
         \pipeline/RegFile_DEC_WB/RegBank[17][0] ,
         \pipeline/RegFile_DEC_WB/RegBank[17][1] ,
         \pipeline/RegFile_DEC_WB/RegBank[17][2] ,
         \pipeline/RegFile_DEC_WB/RegBank[17][3] ,
         \pipeline/RegFile_DEC_WB/RegBank[17][4] ,
         \pipeline/RegFile_DEC_WB/RegBank[17][5] ,
         \pipeline/RegFile_DEC_WB/RegBank[17][6] ,
         \pipeline/RegFile_DEC_WB/RegBank[17][7] ,
         \pipeline/RegFile_DEC_WB/RegBank[17][8] ,
         \pipeline/RegFile_DEC_WB/RegBank[17][9] ,
         \pipeline/RegFile_DEC_WB/RegBank[17][10] ,
         \pipeline/RegFile_DEC_WB/RegBank[17][11] ,
         \pipeline/RegFile_DEC_WB/RegBank[17][12] ,
         \pipeline/RegFile_DEC_WB/RegBank[17][13] ,
         \pipeline/RegFile_DEC_WB/RegBank[17][14] ,
         \pipeline/RegFile_DEC_WB/RegBank[17][15] ,
         \pipeline/RegFile_DEC_WB/RegBank[17][16] ,
         \pipeline/RegFile_DEC_WB/RegBank[17][17] ,
         \pipeline/RegFile_DEC_WB/RegBank[17][18] ,
         \pipeline/RegFile_DEC_WB/RegBank[17][19] ,
         \pipeline/RegFile_DEC_WB/RegBank[17][20] ,
         \pipeline/RegFile_DEC_WB/RegBank[17][21] ,
         \pipeline/RegFile_DEC_WB/RegBank[17][22] ,
         \pipeline/RegFile_DEC_WB/RegBank[17][23] ,
         \pipeline/RegFile_DEC_WB/RegBank[17][24] ,
         \pipeline/RegFile_DEC_WB/RegBank[17][25] ,
         \pipeline/RegFile_DEC_WB/RegBank[17][26] ,
         \pipeline/RegFile_DEC_WB/RegBank[17][27] ,
         \pipeline/RegFile_DEC_WB/RegBank[17][28] ,
         \pipeline/RegFile_DEC_WB/RegBank[17][29] ,
         \pipeline/RegFile_DEC_WB/RegBank[17][30] ,
         \pipeline/RegFile_DEC_WB/RegBank[17][31] ,
         \pipeline/RegFile_DEC_WB/RegBank[16][0] ,
         \pipeline/RegFile_DEC_WB/RegBank[16][1] ,
         \pipeline/RegFile_DEC_WB/RegBank[16][2] ,
         \pipeline/RegFile_DEC_WB/RegBank[16][3] ,
         \pipeline/RegFile_DEC_WB/RegBank[16][4] ,
         \pipeline/RegFile_DEC_WB/RegBank[16][5] ,
         \pipeline/RegFile_DEC_WB/RegBank[16][6] ,
         \pipeline/RegFile_DEC_WB/RegBank[16][7] ,
         \pipeline/RegFile_DEC_WB/RegBank[16][8] ,
         \pipeline/RegFile_DEC_WB/RegBank[16][9] ,
         \pipeline/RegFile_DEC_WB/RegBank[16][10] ,
         \pipeline/RegFile_DEC_WB/RegBank[16][11] ,
         \pipeline/RegFile_DEC_WB/RegBank[16][12] ,
         \pipeline/RegFile_DEC_WB/RegBank[16][13] ,
         \pipeline/RegFile_DEC_WB/RegBank[16][14] ,
         \pipeline/RegFile_DEC_WB/RegBank[16][15] ,
         \pipeline/RegFile_DEC_WB/RegBank[16][16] ,
         \pipeline/RegFile_DEC_WB/RegBank[16][17] ,
         \pipeline/RegFile_DEC_WB/RegBank[16][18] ,
         \pipeline/RegFile_DEC_WB/RegBank[16][19] ,
         \pipeline/RegFile_DEC_WB/RegBank[16][20] ,
         \pipeline/RegFile_DEC_WB/RegBank[16][21] ,
         \pipeline/RegFile_DEC_WB/RegBank[16][22] ,
         \pipeline/RegFile_DEC_WB/RegBank[16][23] ,
         \pipeline/RegFile_DEC_WB/RegBank[16][24] ,
         \pipeline/RegFile_DEC_WB/RegBank[16][25] ,
         \pipeline/RegFile_DEC_WB/RegBank[16][26] ,
         \pipeline/RegFile_DEC_WB/RegBank[16][27] ,
         \pipeline/RegFile_DEC_WB/RegBank[16][28] ,
         \pipeline/RegFile_DEC_WB/RegBank[16][29] ,
         \pipeline/RegFile_DEC_WB/RegBank[16][30] ,
         \pipeline/RegFile_DEC_WB/RegBank[16][31] ,
         \pipeline/RegFile_DEC_WB/RegBank[15][0] ,
         \pipeline/RegFile_DEC_WB/RegBank[15][1] ,
         \pipeline/RegFile_DEC_WB/RegBank[15][2] ,
         \pipeline/RegFile_DEC_WB/RegBank[15][3] ,
         \pipeline/RegFile_DEC_WB/RegBank[15][4] ,
         \pipeline/RegFile_DEC_WB/RegBank[15][5] ,
         \pipeline/RegFile_DEC_WB/RegBank[15][6] ,
         \pipeline/RegFile_DEC_WB/RegBank[15][7] ,
         \pipeline/RegFile_DEC_WB/RegBank[15][8] ,
         \pipeline/RegFile_DEC_WB/RegBank[15][9] ,
         \pipeline/RegFile_DEC_WB/RegBank[15][10] ,
         \pipeline/RegFile_DEC_WB/RegBank[15][11] ,
         \pipeline/RegFile_DEC_WB/RegBank[15][12] ,
         \pipeline/RegFile_DEC_WB/RegBank[15][13] ,
         \pipeline/RegFile_DEC_WB/RegBank[15][14] ,
         \pipeline/RegFile_DEC_WB/RegBank[15][15] ,
         \pipeline/RegFile_DEC_WB/RegBank[15][16] ,
         \pipeline/RegFile_DEC_WB/RegBank[15][17] ,
         \pipeline/RegFile_DEC_WB/RegBank[15][18] ,
         \pipeline/RegFile_DEC_WB/RegBank[15][19] ,
         \pipeline/RegFile_DEC_WB/RegBank[15][20] ,
         \pipeline/RegFile_DEC_WB/RegBank[15][21] ,
         \pipeline/RegFile_DEC_WB/RegBank[15][22] ,
         \pipeline/RegFile_DEC_WB/RegBank[15][23] ,
         \pipeline/RegFile_DEC_WB/RegBank[15][24] ,
         \pipeline/RegFile_DEC_WB/RegBank[15][25] ,
         \pipeline/RegFile_DEC_WB/RegBank[15][26] ,
         \pipeline/RegFile_DEC_WB/RegBank[15][27] ,
         \pipeline/RegFile_DEC_WB/RegBank[15][28] ,
         \pipeline/RegFile_DEC_WB/RegBank[15][29] ,
         \pipeline/RegFile_DEC_WB/RegBank[15][30] ,
         \pipeline/RegFile_DEC_WB/RegBank[15][31] ,
         \pipeline/RegFile_DEC_WB/RegBank[14][0] ,
         \pipeline/RegFile_DEC_WB/RegBank[14][1] ,
         \pipeline/RegFile_DEC_WB/RegBank[14][2] ,
         \pipeline/RegFile_DEC_WB/RegBank[14][3] ,
         \pipeline/RegFile_DEC_WB/RegBank[14][4] ,
         \pipeline/RegFile_DEC_WB/RegBank[14][5] ,
         \pipeline/RegFile_DEC_WB/RegBank[14][6] ,
         \pipeline/RegFile_DEC_WB/RegBank[14][7] ,
         \pipeline/RegFile_DEC_WB/RegBank[14][8] ,
         \pipeline/RegFile_DEC_WB/RegBank[14][9] ,
         \pipeline/RegFile_DEC_WB/RegBank[14][10] ,
         \pipeline/RegFile_DEC_WB/RegBank[14][11] ,
         \pipeline/RegFile_DEC_WB/RegBank[14][12] ,
         \pipeline/RegFile_DEC_WB/RegBank[14][13] ,
         \pipeline/RegFile_DEC_WB/RegBank[14][14] ,
         \pipeline/RegFile_DEC_WB/RegBank[14][15] ,
         \pipeline/RegFile_DEC_WB/RegBank[14][16] ,
         \pipeline/RegFile_DEC_WB/RegBank[14][17] ,
         \pipeline/RegFile_DEC_WB/RegBank[14][18] ,
         \pipeline/RegFile_DEC_WB/RegBank[14][19] ,
         \pipeline/RegFile_DEC_WB/RegBank[14][20] ,
         \pipeline/RegFile_DEC_WB/RegBank[14][21] ,
         \pipeline/RegFile_DEC_WB/RegBank[14][22] ,
         \pipeline/RegFile_DEC_WB/RegBank[14][23] ,
         \pipeline/RegFile_DEC_WB/RegBank[14][24] ,
         \pipeline/RegFile_DEC_WB/RegBank[14][25] ,
         \pipeline/RegFile_DEC_WB/RegBank[14][26] ,
         \pipeline/RegFile_DEC_WB/RegBank[14][27] ,
         \pipeline/RegFile_DEC_WB/RegBank[14][28] ,
         \pipeline/RegFile_DEC_WB/RegBank[14][29] ,
         \pipeline/RegFile_DEC_WB/RegBank[14][30] ,
         \pipeline/RegFile_DEC_WB/RegBank[14][31] ,
         \pipeline/RegFile_DEC_WB/RegBank[13][0] ,
         \pipeline/RegFile_DEC_WB/RegBank[13][1] ,
         \pipeline/RegFile_DEC_WB/RegBank[13][2] ,
         \pipeline/RegFile_DEC_WB/RegBank[13][3] ,
         \pipeline/RegFile_DEC_WB/RegBank[13][4] ,
         \pipeline/RegFile_DEC_WB/RegBank[13][5] ,
         \pipeline/RegFile_DEC_WB/RegBank[13][6] ,
         \pipeline/RegFile_DEC_WB/RegBank[13][7] ,
         \pipeline/RegFile_DEC_WB/RegBank[13][8] ,
         \pipeline/RegFile_DEC_WB/RegBank[13][9] ,
         \pipeline/RegFile_DEC_WB/RegBank[13][10] ,
         \pipeline/RegFile_DEC_WB/RegBank[13][11] ,
         \pipeline/RegFile_DEC_WB/RegBank[13][12] ,
         \pipeline/RegFile_DEC_WB/RegBank[13][13] ,
         \pipeline/RegFile_DEC_WB/RegBank[13][14] ,
         \pipeline/RegFile_DEC_WB/RegBank[13][15] ,
         \pipeline/RegFile_DEC_WB/RegBank[13][16] ,
         \pipeline/RegFile_DEC_WB/RegBank[13][17] ,
         \pipeline/RegFile_DEC_WB/RegBank[13][18] ,
         \pipeline/RegFile_DEC_WB/RegBank[13][19] ,
         \pipeline/RegFile_DEC_WB/RegBank[13][20] ,
         \pipeline/RegFile_DEC_WB/RegBank[13][21] ,
         \pipeline/RegFile_DEC_WB/RegBank[13][22] ,
         \pipeline/RegFile_DEC_WB/RegBank[13][23] ,
         \pipeline/RegFile_DEC_WB/RegBank[13][24] ,
         \pipeline/RegFile_DEC_WB/RegBank[13][25] ,
         \pipeline/RegFile_DEC_WB/RegBank[13][26] ,
         \pipeline/RegFile_DEC_WB/RegBank[13][27] ,
         \pipeline/RegFile_DEC_WB/RegBank[13][28] ,
         \pipeline/RegFile_DEC_WB/RegBank[13][29] ,
         \pipeline/RegFile_DEC_WB/RegBank[13][30] ,
         \pipeline/RegFile_DEC_WB/RegBank[13][31] ,
         \pipeline/RegFile_DEC_WB/RegBank[12][0] ,
         \pipeline/RegFile_DEC_WB/RegBank[12][1] ,
         \pipeline/RegFile_DEC_WB/RegBank[12][2] ,
         \pipeline/RegFile_DEC_WB/RegBank[12][3] ,
         \pipeline/RegFile_DEC_WB/RegBank[12][4] ,
         \pipeline/RegFile_DEC_WB/RegBank[12][5] ,
         \pipeline/RegFile_DEC_WB/RegBank[12][6] ,
         \pipeline/RegFile_DEC_WB/RegBank[12][7] ,
         \pipeline/RegFile_DEC_WB/RegBank[12][8] ,
         \pipeline/RegFile_DEC_WB/RegBank[12][9] ,
         \pipeline/RegFile_DEC_WB/RegBank[12][10] ,
         \pipeline/RegFile_DEC_WB/RegBank[12][11] ,
         \pipeline/RegFile_DEC_WB/RegBank[12][12] ,
         \pipeline/RegFile_DEC_WB/RegBank[12][13] ,
         \pipeline/RegFile_DEC_WB/RegBank[12][14] ,
         \pipeline/RegFile_DEC_WB/RegBank[12][15] ,
         \pipeline/RegFile_DEC_WB/RegBank[12][16] ,
         \pipeline/RegFile_DEC_WB/RegBank[12][17] ,
         \pipeline/RegFile_DEC_WB/RegBank[12][18] ,
         \pipeline/RegFile_DEC_WB/RegBank[12][19] ,
         \pipeline/RegFile_DEC_WB/RegBank[12][20] ,
         \pipeline/RegFile_DEC_WB/RegBank[12][21] ,
         \pipeline/RegFile_DEC_WB/RegBank[12][22] ,
         \pipeline/RegFile_DEC_WB/RegBank[12][23] ,
         \pipeline/RegFile_DEC_WB/RegBank[12][24] ,
         \pipeline/RegFile_DEC_WB/RegBank[12][25] ,
         \pipeline/RegFile_DEC_WB/RegBank[12][26] ,
         \pipeline/RegFile_DEC_WB/RegBank[12][27] ,
         \pipeline/RegFile_DEC_WB/RegBank[12][28] ,
         \pipeline/RegFile_DEC_WB/RegBank[12][29] ,
         \pipeline/RegFile_DEC_WB/RegBank[12][30] ,
         \pipeline/RegFile_DEC_WB/RegBank[12][31] ,
         \pipeline/RegFile_DEC_WB/RegBank[11][0] ,
         \pipeline/RegFile_DEC_WB/RegBank[11][1] ,
         \pipeline/RegFile_DEC_WB/RegBank[11][2] ,
         \pipeline/RegFile_DEC_WB/RegBank[11][3] ,
         \pipeline/RegFile_DEC_WB/RegBank[11][4] ,
         \pipeline/RegFile_DEC_WB/RegBank[11][5] ,
         \pipeline/RegFile_DEC_WB/RegBank[11][6] ,
         \pipeline/RegFile_DEC_WB/RegBank[11][7] ,
         \pipeline/RegFile_DEC_WB/RegBank[11][8] ,
         \pipeline/RegFile_DEC_WB/RegBank[11][9] ,
         \pipeline/RegFile_DEC_WB/RegBank[11][10] ,
         \pipeline/RegFile_DEC_WB/RegBank[11][11] ,
         \pipeline/RegFile_DEC_WB/RegBank[11][12] ,
         \pipeline/RegFile_DEC_WB/RegBank[11][13] ,
         \pipeline/RegFile_DEC_WB/RegBank[11][14] ,
         \pipeline/RegFile_DEC_WB/RegBank[11][15] ,
         \pipeline/RegFile_DEC_WB/RegBank[11][16] ,
         \pipeline/RegFile_DEC_WB/RegBank[11][17] ,
         \pipeline/RegFile_DEC_WB/RegBank[11][18] ,
         \pipeline/RegFile_DEC_WB/RegBank[11][19] ,
         \pipeline/RegFile_DEC_WB/RegBank[11][20] ,
         \pipeline/RegFile_DEC_WB/RegBank[11][21] ,
         \pipeline/RegFile_DEC_WB/RegBank[11][22] ,
         \pipeline/RegFile_DEC_WB/RegBank[11][23] ,
         \pipeline/RegFile_DEC_WB/RegBank[11][24] ,
         \pipeline/RegFile_DEC_WB/RegBank[11][25] ,
         \pipeline/RegFile_DEC_WB/RegBank[11][26] ,
         \pipeline/RegFile_DEC_WB/RegBank[11][27] ,
         \pipeline/RegFile_DEC_WB/RegBank[11][28] ,
         \pipeline/RegFile_DEC_WB/RegBank[11][29] ,
         \pipeline/RegFile_DEC_WB/RegBank[11][30] ,
         \pipeline/RegFile_DEC_WB/RegBank[11][31] ,
         \pipeline/RegFile_DEC_WB/RegBank[10][0] ,
         \pipeline/RegFile_DEC_WB/RegBank[10][1] ,
         \pipeline/RegFile_DEC_WB/RegBank[10][2] ,
         \pipeline/RegFile_DEC_WB/RegBank[10][3] ,
         \pipeline/RegFile_DEC_WB/RegBank[10][4] ,
         \pipeline/RegFile_DEC_WB/RegBank[10][5] ,
         \pipeline/RegFile_DEC_WB/RegBank[10][6] ,
         \pipeline/RegFile_DEC_WB/RegBank[10][7] ,
         \pipeline/RegFile_DEC_WB/RegBank[10][8] ,
         \pipeline/RegFile_DEC_WB/RegBank[10][9] ,
         \pipeline/RegFile_DEC_WB/RegBank[10][10] ,
         \pipeline/RegFile_DEC_WB/RegBank[10][11] ,
         \pipeline/RegFile_DEC_WB/RegBank[10][12] ,
         \pipeline/RegFile_DEC_WB/RegBank[10][13] ,
         \pipeline/RegFile_DEC_WB/RegBank[10][14] ,
         \pipeline/RegFile_DEC_WB/RegBank[10][15] ,
         \pipeline/RegFile_DEC_WB/RegBank[10][16] ,
         \pipeline/RegFile_DEC_WB/RegBank[10][17] ,
         \pipeline/RegFile_DEC_WB/RegBank[10][18] ,
         \pipeline/RegFile_DEC_WB/RegBank[10][19] ,
         \pipeline/RegFile_DEC_WB/RegBank[10][20] ,
         \pipeline/RegFile_DEC_WB/RegBank[10][21] ,
         \pipeline/RegFile_DEC_WB/RegBank[10][22] ,
         \pipeline/RegFile_DEC_WB/RegBank[10][23] ,
         \pipeline/RegFile_DEC_WB/RegBank[10][24] ,
         \pipeline/RegFile_DEC_WB/RegBank[10][25] ,
         \pipeline/RegFile_DEC_WB/RegBank[10][26] ,
         \pipeline/RegFile_DEC_WB/RegBank[10][27] ,
         \pipeline/RegFile_DEC_WB/RegBank[10][28] ,
         \pipeline/RegFile_DEC_WB/RegBank[10][29] ,
         \pipeline/RegFile_DEC_WB/RegBank[10][30] ,
         \pipeline/RegFile_DEC_WB/RegBank[10][31] ,
         \pipeline/RegFile_DEC_WB/RegBank[9][0] ,
         \pipeline/RegFile_DEC_WB/RegBank[9][1] ,
         \pipeline/RegFile_DEC_WB/RegBank[9][2] ,
         \pipeline/RegFile_DEC_WB/RegBank[9][3] ,
         \pipeline/RegFile_DEC_WB/RegBank[9][4] ,
         \pipeline/RegFile_DEC_WB/RegBank[9][5] ,
         \pipeline/RegFile_DEC_WB/RegBank[9][6] ,
         \pipeline/RegFile_DEC_WB/RegBank[9][7] ,
         \pipeline/RegFile_DEC_WB/RegBank[9][8] ,
         \pipeline/RegFile_DEC_WB/RegBank[9][9] ,
         \pipeline/RegFile_DEC_WB/RegBank[9][10] ,
         \pipeline/RegFile_DEC_WB/RegBank[9][11] ,
         \pipeline/RegFile_DEC_WB/RegBank[9][12] ,
         \pipeline/RegFile_DEC_WB/RegBank[9][13] ,
         \pipeline/RegFile_DEC_WB/RegBank[9][14] ,
         \pipeline/RegFile_DEC_WB/RegBank[9][15] ,
         \pipeline/RegFile_DEC_WB/RegBank[9][16] ,
         \pipeline/RegFile_DEC_WB/RegBank[9][17] ,
         \pipeline/RegFile_DEC_WB/RegBank[9][18] ,
         \pipeline/RegFile_DEC_WB/RegBank[9][19] ,
         \pipeline/RegFile_DEC_WB/RegBank[9][20] ,
         \pipeline/RegFile_DEC_WB/RegBank[9][21] ,
         \pipeline/RegFile_DEC_WB/RegBank[9][22] ,
         \pipeline/RegFile_DEC_WB/RegBank[9][23] ,
         \pipeline/RegFile_DEC_WB/RegBank[9][24] ,
         \pipeline/RegFile_DEC_WB/RegBank[9][25] ,
         \pipeline/RegFile_DEC_WB/RegBank[9][26] ,
         \pipeline/RegFile_DEC_WB/RegBank[9][27] ,
         \pipeline/RegFile_DEC_WB/RegBank[9][28] ,
         \pipeline/RegFile_DEC_WB/RegBank[9][29] ,
         \pipeline/RegFile_DEC_WB/RegBank[9][30] ,
         \pipeline/RegFile_DEC_WB/RegBank[9][31] ,
         \pipeline/RegFile_DEC_WB/RegBank[8][0] ,
         \pipeline/RegFile_DEC_WB/RegBank[8][1] ,
         \pipeline/RegFile_DEC_WB/RegBank[8][2] ,
         \pipeline/RegFile_DEC_WB/RegBank[8][3] ,
         \pipeline/RegFile_DEC_WB/RegBank[8][4] ,
         \pipeline/RegFile_DEC_WB/RegBank[8][5] ,
         \pipeline/RegFile_DEC_WB/RegBank[8][6] ,
         \pipeline/RegFile_DEC_WB/RegBank[8][7] ,
         \pipeline/RegFile_DEC_WB/RegBank[8][8] ,
         \pipeline/RegFile_DEC_WB/RegBank[8][9] ,
         \pipeline/RegFile_DEC_WB/RegBank[8][10] ,
         \pipeline/RegFile_DEC_WB/RegBank[8][11] ,
         \pipeline/RegFile_DEC_WB/RegBank[8][12] ,
         \pipeline/RegFile_DEC_WB/RegBank[8][13] ,
         \pipeline/RegFile_DEC_WB/RegBank[8][14] ,
         \pipeline/RegFile_DEC_WB/RegBank[8][15] ,
         \pipeline/RegFile_DEC_WB/RegBank[8][16] ,
         \pipeline/RegFile_DEC_WB/RegBank[8][17] ,
         \pipeline/RegFile_DEC_WB/RegBank[8][18] ,
         \pipeline/RegFile_DEC_WB/RegBank[8][19] ,
         \pipeline/RegFile_DEC_WB/RegBank[8][20] ,
         \pipeline/RegFile_DEC_WB/RegBank[8][21] ,
         \pipeline/RegFile_DEC_WB/RegBank[8][22] ,
         \pipeline/RegFile_DEC_WB/RegBank[8][23] ,
         \pipeline/RegFile_DEC_WB/RegBank[8][24] ,
         \pipeline/RegFile_DEC_WB/RegBank[8][25] ,
         \pipeline/RegFile_DEC_WB/RegBank[8][26] ,
         \pipeline/RegFile_DEC_WB/RegBank[8][27] ,
         \pipeline/RegFile_DEC_WB/RegBank[8][28] ,
         \pipeline/RegFile_DEC_WB/RegBank[8][29] ,
         \pipeline/RegFile_DEC_WB/RegBank[8][30] ,
         \pipeline/RegFile_DEC_WB/RegBank[8][31] ,
         \pipeline/RegFile_DEC_WB/RegBank[7][0] ,
         \pipeline/RegFile_DEC_WB/RegBank[7][1] ,
         \pipeline/RegFile_DEC_WB/RegBank[7][2] ,
         \pipeline/RegFile_DEC_WB/RegBank[7][3] ,
         \pipeline/RegFile_DEC_WB/RegBank[7][4] ,
         \pipeline/RegFile_DEC_WB/RegBank[7][5] ,
         \pipeline/RegFile_DEC_WB/RegBank[7][6] ,
         \pipeline/RegFile_DEC_WB/RegBank[7][7] ,
         \pipeline/RegFile_DEC_WB/RegBank[7][8] ,
         \pipeline/RegFile_DEC_WB/RegBank[7][9] ,
         \pipeline/RegFile_DEC_WB/RegBank[7][10] ,
         \pipeline/RegFile_DEC_WB/RegBank[7][11] ,
         \pipeline/RegFile_DEC_WB/RegBank[7][12] ,
         \pipeline/RegFile_DEC_WB/RegBank[7][13] ,
         \pipeline/RegFile_DEC_WB/RegBank[7][14] ,
         \pipeline/RegFile_DEC_WB/RegBank[7][15] ,
         \pipeline/RegFile_DEC_WB/RegBank[7][16] ,
         \pipeline/RegFile_DEC_WB/RegBank[7][17] ,
         \pipeline/RegFile_DEC_WB/RegBank[7][18] ,
         \pipeline/RegFile_DEC_WB/RegBank[7][19] ,
         \pipeline/RegFile_DEC_WB/RegBank[7][20] ,
         \pipeline/RegFile_DEC_WB/RegBank[7][21] ,
         \pipeline/RegFile_DEC_WB/RegBank[7][22] ,
         \pipeline/RegFile_DEC_WB/RegBank[7][23] ,
         \pipeline/RegFile_DEC_WB/RegBank[7][24] ,
         \pipeline/RegFile_DEC_WB/RegBank[7][25] ,
         \pipeline/RegFile_DEC_WB/RegBank[7][26] ,
         \pipeline/RegFile_DEC_WB/RegBank[7][27] ,
         \pipeline/RegFile_DEC_WB/RegBank[7][28] ,
         \pipeline/RegFile_DEC_WB/RegBank[7][29] ,
         \pipeline/RegFile_DEC_WB/RegBank[7][30] ,
         \pipeline/RegFile_DEC_WB/RegBank[7][31] ,
         \pipeline/RegFile_DEC_WB/RegBank[6][0] ,
         \pipeline/RegFile_DEC_WB/RegBank[6][1] ,
         \pipeline/RegFile_DEC_WB/RegBank[6][2] ,
         \pipeline/RegFile_DEC_WB/RegBank[6][3] ,
         \pipeline/RegFile_DEC_WB/RegBank[6][4] ,
         \pipeline/RegFile_DEC_WB/RegBank[6][5] ,
         \pipeline/RegFile_DEC_WB/RegBank[6][6] ,
         \pipeline/RegFile_DEC_WB/RegBank[6][7] ,
         \pipeline/RegFile_DEC_WB/RegBank[6][8] ,
         \pipeline/RegFile_DEC_WB/RegBank[6][9] ,
         \pipeline/RegFile_DEC_WB/RegBank[6][10] ,
         \pipeline/RegFile_DEC_WB/RegBank[6][11] ,
         \pipeline/RegFile_DEC_WB/RegBank[6][12] ,
         \pipeline/RegFile_DEC_WB/RegBank[6][13] ,
         \pipeline/RegFile_DEC_WB/RegBank[6][14] ,
         \pipeline/RegFile_DEC_WB/RegBank[6][15] ,
         \pipeline/RegFile_DEC_WB/RegBank[6][16] ,
         \pipeline/RegFile_DEC_WB/RegBank[6][17] ,
         \pipeline/RegFile_DEC_WB/RegBank[6][18] ,
         \pipeline/RegFile_DEC_WB/RegBank[6][19] ,
         \pipeline/RegFile_DEC_WB/RegBank[6][20] ,
         \pipeline/RegFile_DEC_WB/RegBank[6][21] ,
         \pipeline/RegFile_DEC_WB/RegBank[6][22] ,
         \pipeline/RegFile_DEC_WB/RegBank[6][23] ,
         \pipeline/RegFile_DEC_WB/RegBank[6][24] ,
         \pipeline/RegFile_DEC_WB/RegBank[6][25] ,
         \pipeline/RegFile_DEC_WB/RegBank[6][26] ,
         \pipeline/RegFile_DEC_WB/RegBank[6][27] ,
         \pipeline/RegFile_DEC_WB/RegBank[6][28] ,
         \pipeline/RegFile_DEC_WB/RegBank[6][29] ,
         \pipeline/RegFile_DEC_WB/RegBank[6][30] ,
         \pipeline/RegFile_DEC_WB/RegBank[6][31] ,
         \pipeline/RegFile_DEC_WB/RegBank[5][0] ,
         \pipeline/RegFile_DEC_WB/RegBank[5][1] ,
         \pipeline/RegFile_DEC_WB/RegBank[5][2] ,
         \pipeline/RegFile_DEC_WB/RegBank[5][3] ,
         \pipeline/RegFile_DEC_WB/RegBank[5][4] ,
         \pipeline/RegFile_DEC_WB/RegBank[5][5] ,
         \pipeline/RegFile_DEC_WB/RegBank[5][6] ,
         \pipeline/RegFile_DEC_WB/RegBank[5][7] ,
         \pipeline/RegFile_DEC_WB/RegBank[5][8] ,
         \pipeline/RegFile_DEC_WB/RegBank[5][9] ,
         \pipeline/RegFile_DEC_WB/RegBank[5][10] ,
         \pipeline/RegFile_DEC_WB/RegBank[5][11] ,
         \pipeline/RegFile_DEC_WB/RegBank[5][12] ,
         \pipeline/RegFile_DEC_WB/RegBank[5][13] ,
         \pipeline/RegFile_DEC_WB/RegBank[5][14] ,
         \pipeline/RegFile_DEC_WB/RegBank[5][15] ,
         \pipeline/RegFile_DEC_WB/RegBank[5][16] ,
         \pipeline/RegFile_DEC_WB/RegBank[5][17] ,
         \pipeline/RegFile_DEC_WB/RegBank[5][18] ,
         \pipeline/RegFile_DEC_WB/RegBank[5][19] ,
         \pipeline/RegFile_DEC_WB/RegBank[5][20] ,
         \pipeline/RegFile_DEC_WB/RegBank[5][21] ,
         \pipeline/RegFile_DEC_WB/RegBank[5][22] ,
         \pipeline/RegFile_DEC_WB/RegBank[5][23] ,
         \pipeline/RegFile_DEC_WB/RegBank[5][24] ,
         \pipeline/RegFile_DEC_WB/RegBank[5][25] ,
         \pipeline/RegFile_DEC_WB/RegBank[5][26] ,
         \pipeline/RegFile_DEC_WB/RegBank[5][27] ,
         \pipeline/RegFile_DEC_WB/RegBank[5][28] ,
         \pipeline/RegFile_DEC_WB/RegBank[5][29] ,
         \pipeline/RegFile_DEC_WB/RegBank[5][30] ,
         \pipeline/RegFile_DEC_WB/RegBank[5][31] ,
         \pipeline/RegFile_DEC_WB/RegBank[4][0] ,
         \pipeline/RegFile_DEC_WB/RegBank[4][1] ,
         \pipeline/RegFile_DEC_WB/RegBank[4][2] ,
         \pipeline/RegFile_DEC_WB/RegBank[4][3] ,
         \pipeline/RegFile_DEC_WB/RegBank[4][4] ,
         \pipeline/RegFile_DEC_WB/RegBank[4][5] ,
         \pipeline/RegFile_DEC_WB/RegBank[4][6] ,
         \pipeline/RegFile_DEC_WB/RegBank[4][7] ,
         \pipeline/RegFile_DEC_WB/RegBank[4][8] ,
         \pipeline/RegFile_DEC_WB/RegBank[4][9] ,
         \pipeline/RegFile_DEC_WB/RegBank[4][10] ,
         \pipeline/RegFile_DEC_WB/RegBank[4][11] ,
         \pipeline/RegFile_DEC_WB/RegBank[4][12] ,
         \pipeline/RegFile_DEC_WB/RegBank[4][13] ,
         \pipeline/RegFile_DEC_WB/RegBank[4][14] ,
         \pipeline/RegFile_DEC_WB/RegBank[4][15] ,
         \pipeline/RegFile_DEC_WB/RegBank[4][16] ,
         \pipeline/RegFile_DEC_WB/RegBank[4][17] ,
         \pipeline/RegFile_DEC_WB/RegBank[4][18] ,
         \pipeline/RegFile_DEC_WB/RegBank[4][19] ,
         \pipeline/RegFile_DEC_WB/RegBank[4][20] ,
         \pipeline/RegFile_DEC_WB/RegBank[4][21] ,
         \pipeline/RegFile_DEC_WB/RegBank[4][22] ,
         \pipeline/RegFile_DEC_WB/RegBank[4][23] ,
         \pipeline/RegFile_DEC_WB/RegBank[4][24] ,
         \pipeline/RegFile_DEC_WB/RegBank[4][25] ,
         \pipeline/RegFile_DEC_WB/RegBank[4][26] ,
         \pipeline/RegFile_DEC_WB/RegBank[4][27] ,
         \pipeline/RegFile_DEC_WB/RegBank[4][28] ,
         \pipeline/RegFile_DEC_WB/RegBank[4][29] ,
         \pipeline/RegFile_DEC_WB/RegBank[4][30] ,
         \pipeline/RegFile_DEC_WB/RegBank[4][31] ,
         \pipeline/RegFile_DEC_WB/RegBank[3][0] ,
         \pipeline/RegFile_DEC_WB/RegBank[3][1] ,
         \pipeline/RegFile_DEC_WB/RegBank[3][2] ,
         \pipeline/RegFile_DEC_WB/RegBank[3][3] ,
         \pipeline/RegFile_DEC_WB/RegBank[3][4] ,
         \pipeline/RegFile_DEC_WB/RegBank[3][5] ,
         \pipeline/RegFile_DEC_WB/RegBank[3][6] ,
         \pipeline/RegFile_DEC_WB/RegBank[3][7] ,
         \pipeline/RegFile_DEC_WB/RegBank[3][8] ,
         \pipeline/RegFile_DEC_WB/RegBank[3][9] ,
         \pipeline/RegFile_DEC_WB/RegBank[3][10] ,
         \pipeline/RegFile_DEC_WB/RegBank[3][11] ,
         \pipeline/RegFile_DEC_WB/RegBank[3][12] ,
         \pipeline/RegFile_DEC_WB/RegBank[3][13] ,
         \pipeline/RegFile_DEC_WB/RegBank[3][14] ,
         \pipeline/RegFile_DEC_WB/RegBank[3][15] ,
         \pipeline/RegFile_DEC_WB/RegBank[3][16] ,
         \pipeline/RegFile_DEC_WB/RegBank[3][17] ,
         \pipeline/RegFile_DEC_WB/RegBank[3][18] ,
         \pipeline/RegFile_DEC_WB/RegBank[3][19] ,
         \pipeline/RegFile_DEC_WB/RegBank[3][20] ,
         \pipeline/RegFile_DEC_WB/RegBank[3][21] ,
         \pipeline/RegFile_DEC_WB/RegBank[3][22] ,
         \pipeline/RegFile_DEC_WB/RegBank[3][23] ,
         \pipeline/RegFile_DEC_WB/RegBank[3][24] ,
         \pipeline/RegFile_DEC_WB/RegBank[3][25] ,
         \pipeline/RegFile_DEC_WB/RegBank[3][26] ,
         \pipeline/RegFile_DEC_WB/RegBank[3][27] ,
         \pipeline/RegFile_DEC_WB/RegBank[3][28] ,
         \pipeline/RegFile_DEC_WB/RegBank[3][29] ,
         \pipeline/RegFile_DEC_WB/RegBank[3][30] ,
         \pipeline/RegFile_DEC_WB/RegBank[3][31] ,
         \pipeline/RegFile_DEC_WB/RegBank[2][0] ,
         \pipeline/RegFile_DEC_WB/RegBank[2][1] ,
         \pipeline/RegFile_DEC_WB/RegBank[2][2] ,
         \pipeline/RegFile_DEC_WB/RegBank[2][3] ,
         \pipeline/RegFile_DEC_WB/RegBank[2][4] ,
         \pipeline/RegFile_DEC_WB/RegBank[2][5] ,
         \pipeline/RegFile_DEC_WB/RegBank[2][6] ,
         \pipeline/RegFile_DEC_WB/RegBank[2][7] ,
         \pipeline/RegFile_DEC_WB/RegBank[2][8] ,
         \pipeline/RegFile_DEC_WB/RegBank[2][9] ,
         \pipeline/RegFile_DEC_WB/RegBank[2][10] ,
         \pipeline/RegFile_DEC_WB/RegBank[2][11] ,
         \pipeline/RegFile_DEC_WB/RegBank[2][12] ,
         \pipeline/RegFile_DEC_WB/RegBank[2][13] ,
         \pipeline/RegFile_DEC_WB/RegBank[2][14] ,
         \pipeline/RegFile_DEC_WB/RegBank[2][15] ,
         \pipeline/RegFile_DEC_WB/RegBank[2][16] ,
         \pipeline/RegFile_DEC_WB/RegBank[2][17] ,
         \pipeline/RegFile_DEC_WB/RegBank[2][18] ,
         \pipeline/RegFile_DEC_WB/RegBank[2][19] ,
         \pipeline/RegFile_DEC_WB/RegBank[2][20] ,
         \pipeline/RegFile_DEC_WB/RegBank[2][21] ,
         \pipeline/RegFile_DEC_WB/RegBank[2][22] ,
         \pipeline/RegFile_DEC_WB/RegBank[2][23] ,
         \pipeline/RegFile_DEC_WB/RegBank[2][24] ,
         \pipeline/RegFile_DEC_WB/RegBank[2][25] ,
         \pipeline/RegFile_DEC_WB/RegBank[2][26] ,
         \pipeline/RegFile_DEC_WB/RegBank[2][27] ,
         \pipeline/RegFile_DEC_WB/RegBank[2][28] ,
         \pipeline/RegFile_DEC_WB/RegBank[2][29] ,
         \pipeline/RegFile_DEC_WB/RegBank[2][30] ,
         \pipeline/RegFile_DEC_WB/RegBank[2][31] ,
         \pipeline/RegFile_DEC_WB/RegBank[1][0] ,
         \pipeline/RegFile_DEC_WB/RegBank[1][1] ,
         \pipeline/RegFile_DEC_WB/RegBank[1][2] ,
         \pipeline/RegFile_DEC_WB/RegBank[1][3] ,
         \pipeline/RegFile_DEC_WB/RegBank[1][4] ,
         \pipeline/RegFile_DEC_WB/RegBank[1][5] ,
         \pipeline/RegFile_DEC_WB/RegBank[1][6] ,
         \pipeline/RegFile_DEC_WB/RegBank[1][7] ,
         \pipeline/RegFile_DEC_WB/RegBank[1][8] ,
         \pipeline/RegFile_DEC_WB/RegBank[1][9] ,
         \pipeline/RegFile_DEC_WB/RegBank[1][10] ,
         \pipeline/RegFile_DEC_WB/RegBank[1][11] ,
         \pipeline/RegFile_DEC_WB/RegBank[1][12] ,
         \pipeline/RegFile_DEC_WB/RegBank[1][13] ,
         \pipeline/RegFile_DEC_WB/RegBank[1][14] ,
         \pipeline/RegFile_DEC_WB/RegBank[1][15] ,
         \pipeline/RegFile_DEC_WB/RegBank[1][16] ,
         \pipeline/RegFile_DEC_WB/RegBank[1][17] ,
         \pipeline/RegFile_DEC_WB/RegBank[1][18] ,
         \pipeline/RegFile_DEC_WB/RegBank[1][19] ,
         \pipeline/RegFile_DEC_WB/RegBank[1][20] ,
         \pipeline/RegFile_DEC_WB/RegBank[1][21] ,
         \pipeline/RegFile_DEC_WB/RegBank[1][22] ,
         \pipeline/RegFile_DEC_WB/RegBank[1][23] ,
         \pipeline/RegFile_DEC_WB/RegBank[1][24] ,
         \pipeline/RegFile_DEC_WB/RegBank[1][25] ,
         \pipeline/RegFile_DEC_WB/RegBank[1][26] ,
         \pipeline/RegFile_DEC_WB/RegBank[1][27] ,
         \pipeline/RegFile_DEC_WB/RegBank[1][28] ,
         \pipeline/RegFile_DEC_WB/RegBank[1][29] ,
         \pipeline/RegFile_DEC_WB/RegBank[1][30] ,
         \pipeline/RegFile_DEC_WB/RegBank[1][31] , \pipeline/IDEX_Stage/N217 ,
         \pipeline/IDEX_Stage/N216 , \pipeline/IDEX_Stage/N215 ,
         \pipeline/IDEX_Stage/N214 , \pipeline/IDEX_Stage/N213 ,
         \pipeline/IDEX_Stage/N212 , \pipeline/IDEX_Stage/N211 ,
         \pipeline/IDEX_Stage/N210 , \pipeline/IDEX_Stage/N209 ,
         \pipeline/IDEX_Stage/N208 , \pipeline/IDEX_Stage/N207 ,
         \pipeline/IDEX_Stage/N206 , \pipeline/IDEX_Stage/N205 ,
         \pipeline/IDEX_Stage/N204 , \pipeline/IDEX_Stage/N203 ,
         \pipeline/IDEX_Stage/N202 , \pipeline/IDEX_Stage/N201 ,
         \pipeline/IDEX_Stage/N200 , \pipeline/IDEX_Stage/N199 ,
         \pipeline/IDEX_Stage/N198 , \pipeline/IDEX_Stage/N197 ,
         \pipeline/IDEX_Stage/N181 , \pipeline/IDEX_Stage/N180 ,
         \pipeline/IDEX_Stage/N179 , \pipeline/IDEX_Stage/N178 ,
         \pipeline/IDEX_Stage/N177 , \pipeline/IDEX_Stage/N176 ,
         \pipeline/IDEX_Stage/N175 , \pipeline/IDEX_Stage/N174 ,
         \pipeline/IDEX_Stage/N173 , \pipeline/IDEX_Stage/N172 ,
         \pipeline/IDEX_Stage/N171 , \pipeline/IDEX_Stage/N170 ,
         \pipeline/IDEX_Stage/N169 , \pipeline/IDEX_Stage/N168 ,
         \pipeline/IDEX_Stage/N167 , \pipeline/IDEX_Stage/N166 ,
         \pipeline/IDEX_Stage/N165 , \pipeline/IDEX_Stage/N164 ,
         \pipeline/IDEX_Stage/N163 , \pipeline/IDEX_Stage/N162 ,
         \pipeline/IDEX_Stage/N161 , \pipeline/IDEX_Stage/N160 ,
         \pipeline/IDEX_Stage/N159 , \pipeline/IDEX_Stage/N158 ,
         \pipeline/IDEX_Stage/N157 , \pipeline/IDEX_Stage/N156 ,
         \pipeline/IDEX_Stage/N155 , \pipeline/IDEX_Stage/N154 ,
         \pipeline/IDEX_Stage/N153 , \pipeline/IDEX_Stage/N152 ,
         \pipeline/IDEX_Stage/N151 , \pipeline/IDEX_Stage/N150 ,
         \pipeline/IDEX_Stage/N149 , \pipeline/IDEX_Stage/N148 ,
         \pipeline/IDEX_Stage/N147 , \pipeline/IDEX_Stage/N146 ,
         \pipeline/IDEX_Stage/N145 , \pipeline/IDEX_Stage/N144 ,
         \pipeline/IDEX_Stage/N143 , \pipeline/IDEX_Stage/N142 ,
         \pipeline/IDEX_Stage/N141 , \pipeline/IDEX_Stage/N140 ,
         \pipeline/IDEX_Stage/N139 , \pipeline/IDEX_Stage/N138 ,
         \pipeline/IDEX_Stage/N137 , \pipeline/IDEX_Stage/N136 ,
         \pipeline/IDEX_Stage/N135 , \pipeline/IDEX_Stage/N134 ,
         \pipeline/IDEX_Stage/N133 , \pipeline/IDEX_Stage/N132 ,
         \pipeline/IDEX_Stage/N131 , \pipeline/IDEX_Stage/N130 ,
         \pipeline/IDEX_Stage/N129 , \pipeline/IDEX_Stage/N128 ,
         \pipeline/IDEX_Stage/N127 , \pipeline/IDEX_Stage/N126 ,
         \pipeline/IDEX_Stage/N125 , \pipeline/IDEX_Stage/N124 ,
         \pipeline/IDEX_Stage/N123 , \pipeline/IDEX_Stage/N122 ,
         \pipeline/IDEX_Stage/N121 , \pipeline/IDEX_Stage/N120 ,
         \pipeline/IDEX_Stage/N119 , \pipeline/IDEX_Stage/N118 ,
         \pipeline/IDEX_Stage/N117 , \pipeline/IDEX_Stage/N116 ,
         \pipeline/IDEX_Stage/N115 , \pipeline/IDEX_Stage/N114 ,
         \pipeline/IDEX_Stage/N113 , \pipeline/IDEX_Stage/N112 ,
         \pipeline/IDEX_Stage/N111 , \pipeline/IDEX_Stage/N110 ,
         \pipeline/IDEX_Stage/N109 , \pipeline/IDEX_Stage/N108 ,
         \pipeline/IDEX_Stage/N107 , \pipeline/IDEX_Stage/N106 ,
         \pipeline/IDEX_Stage/N105 , \pipeline/IDEX_Stage/N104 ,
         \pipeline/IDEX_Stage/N103 , \pipeline/IDEX_Stage/N102 ,
         \pipeline/IDEX_Stage/N101 , \pipeline/IDEX_Stage/N100 ,
         \pipeline/IDEX_Stage/N99 , \pipeline/IDEX_Stage/N98 ,
         \pipeline/IDEX_Stage/N97 , \pipeline/IDEX_Stage/N96 ,
         \pipeline/IDEX_Stage/N95 , \pipeline/IDEX_Stage/N94 ,
         \pipeline/IDEX_Stage/N93 , \pipeline/IDEX_Stage/N92 ,
         \pipeline/IDEX_Stage/N91 , \pipeline/IDEX_Stage/N90 ,
         \pipeline/IDEX_Stage/N89 , \pipeline/stageE/input2_to_ALU[0] ,
         \pipeline/stageE/EXE_ALU/add_alu/sCout[0] ,
         \pipeline/stageE/EXE_ALU/alu_shift/N265 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N264 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N263 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N262 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N261 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N260 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N259 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N258 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N257 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N256 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N255 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N254 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N253 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N252 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N251 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N250 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N249 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N248 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N247 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N246 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N245 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N244 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N243 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N242 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N241 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N240 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N239 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N238 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N237 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N236 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N235 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N234 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N233 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N232 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N231 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N230 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N229 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N228 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N227 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N226 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N225 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N224 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N223 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N222 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N221 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N220 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N219 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N218 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N217 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N216 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N215 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N214 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N213 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N212 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N211 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N210 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N209 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N208 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N207 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N206 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N205 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N204 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N203 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N202 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N168 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N167 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N166 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N165 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N164 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N163 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N162 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N161 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N160 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N159 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N158 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N157 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N156 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N155 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N154 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N153 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N152 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N151 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N150 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N149 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N148 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N147 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N146 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N145 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N144 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N143 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N142 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N141 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N140 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N139 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N138 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N137 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N136 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N135 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N134 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N133 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N132 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N131 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N130 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N129 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N128 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N127 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N126 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N125 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N124 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N123 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N122 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N121 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N120 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N119 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N118 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N117 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N116 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N115 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N114 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N113 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N112 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N111 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N110 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N109 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N108 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N107 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N106 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N105 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N70 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N69 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N68 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N67 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N66 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N65 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N64 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N63 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N62 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N61 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N60 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N59 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N58 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N57 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N56 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N55 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N54 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N53 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N52 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N51 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N50 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N49 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N48 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N47 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N46 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N45 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N44 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N43 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N42 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N41 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N40 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N39 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N38 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N37 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N36 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N35 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N34 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N33 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N32 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N31 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N30 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N29 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N28 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N27 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N26 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N25 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N24 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N23 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N22 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N21 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N20 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N19 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N18 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N17 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N16 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N15 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N14 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N13 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N12 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N11 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N10 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N9 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N8 ,
         \pipeline/stageE/EXE_ALU/alu_shift/N7 , \pipeline/EXMEM_stage/N76 ,
         \pipeline/EXMEM_stage/N75 , \pipeline/EXMEM_stage/N74 ,
         \pipeline/EXMEM_stage/N73 , \pipeline/EXMEM_stage/N72 ,
         \pipeline/EXMEM_stage/N71 , \pipeline/EXMEM_stage/N70 ,
         \pipeline/EXMEM_stage/N69 , \pipeline/EXMEM_stage/N68 ,
         \pipeline/EXMEM_stage/N67 , \pipeline/EXMEM_stage/N66 ,
         \pipeline/EXMEM_stage/N65 , \pipeline/EXMEM_stage/N64 ,
         \pipeline/EXMEM_stage/N63 , \pipeline/EXMEM_stage/N62 ,
         \pipeline/EXMEM_stage/N61 , \pipeline/EXMEM_stage/N60 ,
         \pipeline/EXMEM_stage/N59 , \pipeline/EXMEM_stage/N58 ,
         \pipeline/EXMEM_stage/N57 , \pipeline/EXMEM_stage/N56 ,
         \pipeline/EXMEM_stage/N55 , \pipeline/EXMEM_stage/N54 ,
         \pipeline/EXMEM_stage/N53 , \pipeline/EXMEM_stage/N52 ,
         \pipeline/EXMEM_stage/N51 , \pipeline/EXMEM_stage/N50 ,
         \pipeline/EXMEM_stage/N49 , \pipeline/EXMEM_stage/N48 ,
         \pipeline/EXMEM_stage/N47 , \pipeline/EXMEM_stage/N46 ,
         \pipeline/EXMEM_stage/N45 , \pipeline/EXMEM_stage/N44 ,
         \pipeline/EXMEM_stage/N43 , \pipeline/EXMEM_stage/N42 ,
         \pipeline/EXMEM_stage/N41 , \pipeline/EXMEM_stage/N40 ,
         \pipeline/EXMEM_stage/N39 , \pipeline/EXMEM_stage/N38 ,
         \pipeline/EXMEM_stage/N37 , \pipeline/EXMEM_stage/N36 ,
         \pipeline/EXMEM_stage/N35 , \pipeline/EXMEM_stage/N34 ,
         \pipeline/EXMEM_stage/N33 , \pipeline/EXMEM_stage/N32 ,
         \pipeline/EXMEM_stage/N31 , \pipeline/EXMEM_stage/N30 ,
         \pipeline/EXMEM_stage/N29 , \pipeline/EXMEM_stage/N28 ,
         \pipeline/EXMEM_stage/N27 , \pipeline/EXMEM_stage/N26 ,
         \pipeline/EXMEM_stage/N25 , \pipeline/EXMEM_stage/N24 ,
         \pipeline/EXMEM_stage/N23 , \pipeline/EXMEM_stage/N22 ,
         \pipeline/EXMEM_stage/N21 , \pipeline/EXMEM_stage/N20 ,
         \pipeline/EXMEM_stage/N19 , \pipeline/EXMEM_stage/N18 ,
         \pipeline/EXMEM_stage/N17 , \pipeline/EXMEM_stage/N16 ,
         \pipeline/EXMEM_stage/N15 , \pipeline/EXMEM_stage/N14 ,
         \pipeline/EXMEM_stage/N13 , \pipeline/EXMEM_stage/N12 ,
         \pipeline/EXMEM_stage/N11 , \pipeline/EXMEM_stage/N10 ,
         \pipeline/EXMEM_stage/N9 , \pipeline/EXMEM_stage/N8 ,
         \pipeline/EXMEM_stage/N7 , \pipeline/EXMEM_stage/N6 ,
         \pipeline/EXMEM_stage/N5 , \pipeline/EXMEM_stage/N4 ,
         \pipeline/EXMEM_stage/N3 , \pipeline/MEMWB_Stage/N47 ,
         \pipeline/MEMWB_Stage/N46 , \pipeline/MEMWB_Stage/N45 ,
         \pipeline/MEMWB_Stage/N44 , \pipeline/MEMWB_Stage/N43 ,
         \pipeline/MEMWB_Stage/N42 , \pipeline/MEMWB_Stage/N41 ,
         \pipeline/MEMWB_Stage/N40 , \pipeline/MEMWB_Stage/N39 ,
         \pipeline/MEMWB_Stage/N38 , \pipeline/MEMWB_Stage/N37 ,
         \pipeline/MEMWB_Stage/N36 , \pipeline/MEMWB_Stage/N35 ,
         \pipeline/MEMWB_Stage/N34 , \pipeline/MEMWB_Stage/N33 ,
         \pipeline/MEMWB_Stage/N32 , \pipeline/MEMWB_Stage/N31 ,
         \pipeline/MEMWB_Stage/N30 , \pipeline/MEMWB_Stage/N29 ,
         \pipeline/MEMWB_Stage/N28 , \pipeline/MEMWB_Stage/N27 ,
         \pipeline/MEMWB_Stage/N26 , \pipeline/MEMWB_Stage/N25 ,
         \pipeline/MEMWB_Stage/N24 , \pipeline/MEMWB_Stage/N23 ,
         \pipeline/MEMWB_Stage/N22 , \pipeline/MEMWB_Stage/N21 ,
         \pipeline/MEMWB_Stage/N20 , \pipeline/MEMWB_Stage/N19 ,
         \pipeline/MEMWB_Stage/N18 , \pipeline/MEMWB_Stage/N17 ,
         \pipeline/MEMWB_Stage/N16 , \pipeline/MEMWB_Stage/N15 ,
         \pipeline/MEMWB_Stage/N14 , \pipeline/MEMWB_Stage/N13 ,
         \pipeline/MEMWB_Stage/N12 , \pipeline/MEMWB_Stage/N11 ,
         \pipeline/MEMWB_Stage/N10 , \pipeline/cu_hazard/N40 ,
         \pipeline/cu_hazard/N39 , \pipeline/cu_pipeline/N113 ,
         \pipeline/cu_pipeline/N112 , \pipeline/cu_pipeline/N110 ,
         \pipeline/cu_pipeline/N109 , \pipeline/cu_pipeline/N108 ,
         \pipeline/cu_pipeline/N107 , \pipeline/cu_pipeline/N106 ,
         \pipeline/cu_pipeline/N105 , \pipeline/cu_pipeline/N104 ,
         \pipeline/cu_pipeline/N103 , \pipeline/cu_pipeline/N102 ,
         \pipeline/cu_pipeline/N101 , \pipeline/cu_pipeline/N89 ,
         \pipeline/cu_pipeline/N88 , \DataMem/N2349 , \DataMem/N2346 ,
         \DataMem/N2343 , \DataMem/N2340 , \DataMem/N2337 , \DataMem/N2334 ,
         \DataMem/N2331 , \DataMem/N2328 , \DataMem/N2325 , \DataMem/N2322 ,
         \DataMem/N2319 , \DataMem/N2316 , \DataMem/N2313 , \DataMem/N2310 ,
         \DataMem/N2307 , \DataMem/N2304 , \DataMem/N2301 , \DataMem/N2298 ,
         \DataMem/N2295 , \DataMem/N2292 , \DataMem/N2289 , \DataMem/N2286 ,
         \DataMem/N2283 , \DataMem/N2280 , \DataMem/N2277 , \DataMem/N2274 ,
         \DataMem/N2271 , \DataMem/N2268 , \DataMem/N2265 , \DataMem/N2262 ,
         \DataMem/N2259 , \DataMem/N2256 , \DataMem/N2254 , \DataMem/N2251 ,
         \DataMem/N2248 , \DataMem/N2245 , \DataMem/N2242 , \DataMem/N2239 ,
         \DataMem/N2236 , \DataMem/N2233 , \DataMem/N2230 , \DataMem/N2227 ,
         \DataMem/N2224 , \DataMem/N2221 , \DataMem/N2218 , \DataMem/N2215 ,
         \DataMem/N2212 , \DataMem/N2209 , \DataMem/N2206 , \DataMem/N2203 ,
         \DataMem/N2200 , \DataMem/N2197 , \DataMem/N2194 , \DataMem/N2191 ,
         \DataMem/N2188 , \DataMem/N2185 , \DataMem/N2182 , \DataMem/N2179 ,
         \DataMem/N2176 , \DataMem/N2173 , \DataMem/N2170 , \DataMem/N2167 ,
         \DataMem/N2164 , \DataMem/N2161 , \DataMem/N2159 , \DataMem/N2157 ,
         \DataMem/N2155 , \DataMem/N2153 , \DataMem/N2151 , \DataMem/N2149 ,
         \DataMem/N2147 , \DataMem/N2145 , \DataMem/N2143 , \DataMem/N2141 ,
         \DataMem/N2139 , \DataMem/N2137 , \DataMem/N2135 , \DataMem/N2133 ,
         \DataMem/N2131 , \DataMem/N2129 , \DataMem/N2127 , \DataMem/N2125 ,
         \DataMem/N2123 , \DataMem/N2121 , \DataMem/N2119 , \DataMem/N2117 ,
         \DataMem/N2115 , \DataMem/N2113 , \DataMem/N2111 , \DataMem/N2109 ,
         \DataMem/N2107 , \DataMem/N2105 , \DataMem/N2103 , \DataMem/N2101 ,
         \DataMem/N2099 , \DataMem/N2097 , \DataMem/N2095 , \DataMem/N2093 ,
         \DataMem/N2091 , \DataMem/N2089 , \DataMem/N2087 , \DataMem/N2085 ,
         \DataMem/N2083 , \DataMem/N2081 , \DataMem/N2079 , \DataMem/N2077 ,
         \DataMem/N2075 , \DataMem/N2073 , \DataMem/N2071 , \DataMem/N2069 ,
         \DataMem/N2067 , \DataMem/N2065 , \DataMem/N2063 , \DataMem/N2061 ,
         \DataMem/N2059 , \DataMem/N2057 , \DataMem/N2055 , \DataMem/N2053 ,
         \DataMem/N2051 , \DataMem/N2049 , \DataMem/N2047 , \DataMem/N2045 ,
         \DataMem/N2043 , \DataMem/N2041 , \DataMem/N2039 , \DataMem/N2037 ,
         \DataMem/N2035 , \DataMem/N2033 , \DataMem/N2031 , \DataMem/N2029 ,
         \DataMem/N2027 , \DataMem/N2025 , \DataMem/N2023 , \DataMem/N2021 ,
         \DataMem/N2019 , \DataMem/N2017 , \DataMem/N2015 , \DataMem/N2013 ,
         \DataMem/N2011 , \DataMem/N2009 , \DataMem/N2007 , \DataMem/N2005 ,
         \DataMem/N2003 , \DataMem/N2001 , \DataMem/N1999 , \DataMem/N1997 ,
         \DataMem/N1995 , \DataMem/N1993 , \DataMem/N1991 , \DataMem/N1989 ,
         \DataMem/N1987 , \DataMem/N1985 , \DataMem/N1983 , \DataMem/N1981 ,
         \DataMem/N1979 , \DataMem/N1977 , \DataMem/N1975 , \DataMem/N1973 ,
         \DataMem/N1971 , \DataMem/N1969 , \DataMem/N1967 , \DataMem/N1965 ,
         \DataMem/N1963 , \DataMem/N1961 , \DataMem/N1959 , \DataMem/N1957 ,
         \DataMem/N1955 , \DataMem/N1953 , \DataMem/N1951 , \DataMem/N1949 ,
         \DataMem/N1947 , \DataMem/N1945 , \DataMem/N1943 , \DataMem/N1941 ,
         \DataMem/N1939 , \DataMem/N1937 , \DataMem/N1935 , \DataMem/N1933 ,
         \DataMem/N1931 , \DataMem/N1929 , \DataMem/N1927 , \DataMem/N1925 ,
         \DataMem/N1923 , \DataMem/N1921 , \DataMem/N1919 , \DataMem/N1917 ,
         \DataMem/N1915 , \DataMem/N1913 , \DataMem/N1911 , \DataMem/N1909 ,
         \DataMem/N1907 , \DataMem/N1905 , \DataMem/N1903 , \DataMem/N1901 ,
         \DataMem/N1899 , \DataMem/N1897 , \DataMem/N1895 , \DataMem/N1893 ,
         \DataMem/N1891 , \DataMem/N1889 , \DataMem/N1887 , \DataMem/N1885 ,
         \DataMem/N1883 , \DataMem/N1881 , \DataMem/N1879 , \DataMem/N1877 ,
         \DataMem/N1875 , \DataMem/N1873 , \DataMem/N1871 , \DataMem/N1869 ,
         \DataMem/N1867 , \DataMem/N1865 , \DataMem/N1863 , \DataMem/N1861 ,
         \DataMem/N1859 , \DataMem/N1857 , \DataMem/N1855 , \DataMem/N1853 ,
         \DataMem/N1851 , \DataMem/N1849 , \DataMem/N1847 , \DataMem/N1845 ,
         \DataMem/N1843 , \DataMem/N1841 , \DataMem/N1839 , \DataMem/N1837 ,
         \DataMem/N1835 , \DataMem/N1833 , \DataMem/N1831 , \DataMem/N1829 ,
         \DataMem/N1827 , \DataMem/N1825 , \DataMem/N1823 , \DataMem/N1821 ,
         \DataMem/N1819 , \DataMem/N1817 , \DataMem/N1815 , \DataMem/N1813 ,
         \DataMem/N1811 , \DataMem/N1809 , \DataMem/N1807 , \DataMem/N1805 ,
         \DataMem/N1803 , \DataMem/N1801 , \DataMem/N1799 , \DataMem/N1797 ,
         \DataMem/N1795 , \DataMem/N1793 , \DataMem/N1791 , \DataMem/N1789 ,
         \DataMem/N1787 , \DataMem/N1785 , \DataMem/N1783 , \DataMem/N1781 ,
         \DataMem/N1779 , \DataMem/N1777 , \DataMem/N1775 , \DataMem/N1773 ,
         \DataMem/N1771 , \DataMem/N1769 , \DataMem/N1767 , \DataMem/N1765 ,
         \DataMem/N1763 , \DataMem/N1761 , \DataMem/N1759 , \DataMem/N1757 ,
         \DataMem/N1755 , \DataMem/N1753 , \DataMem/N1751 , \DataMem/N1749 ,
         \DataMem/N1747 , \DataMem/N1745 , \DataMem/N1743 , \DataMem/N1741 ,
         \DataMem/N1739 , \DataMem/N1737 , \DataMem/N1735 , \DataMem/N1733 ,
         \DataMem/N1731 , \DataMem/N1729 , \DataMem/N1727 , \DataMem/N1725 ,
         \DataMem/N1723 , \DataMem/N1721 , \DataMem/N1719 , \DataMem/N1717 ,
         \DataMem/N1715 , \DataMem/N1713 , \DataMem/N1711 , \DataMem/N1709 ,
         \DataMem/N1707 , \DataMem/N1705 , \DataMem/N1703 , \DataMem/N1701 ,
         \DataMem/N1699 , \DataMem/N1697 , \DataMem/N1695 , \DataMem/N1693 ,
         \DataMem/N1691 , \DataMem/N1689 , \DataMem/N1687 , \DataMem/N1685 ,
         \DataMem/N1683 , \DataMem/N1681 , \DataMem/N1679 , \DataMem/N1677 ,
         \DataMem/N1675 , \DataMem/N1673 , \DataMem/N1671 , \DataMem/N1669 ,
         \DataMem/N1667 , \DataMem/N1665 , \DataMem/N1663 , \DataMem/N1661 ,
         \DataMem/N1659 , \DataMem/N1657 , \DataMem/N1655 , \DataMem/N1653 ,
         \DataMem/N1651 , \DataMem/N1649 , \DataMem/Mem[0][0] ,
         \DataMem/Mem[0][1] , \DataMem/Mem[0][2] , \DataMem/Mem[0][3] ,
         \DataMem/Mem[0][4] , \DataMem/Mem[0][5] , \DataMem/Mem[0][6] ,
         \DataMem/Mem[0][7] , \DataMem/Mem[0][8] , \DataMem/Mem[0][9] ,
         \DataMem/Mem[0][10] , \DataMem/Mem[0][11] , \DataMem/Mem[0][12] ,
         \DataMem/Mem[0][13] , \DataMem/Mem[0][14] , \DataMem/Mem[0][15] ,
         \DataMem/Mem[0][16] , \DataMem/Mem[0][17] , \DataMem/Mem[0][18] ,
         \DataMem/Mem[0][19] , \DataMem/Mem[0][20] , \DataMem/Mem[0][21] ,
         \DataMem/Mem[0][22] , \DataMem/Mem[0][23] , \DataMem/Mem[0][24] ,
         \DataMem/Mem[0][25] , \DataMem/Mem[0][26] , \DataMem/Mem[0][27] ,
         \DataMem/Mem[0][28] , \DataMem/Mem[0][29] , \DataMem/Mem[0][30] ,
         \DataMem/Mem[0][31] , \DataMem/Mem[1][0] , \DataMem/Mem[1][1] ,
         \DataMem/Mem[1][2] , \DataMem/Mem[1][3] , \DataMem/Mem[1][4] ,
         \DataMem/Mem[1][5] , \DataMem/Mem[1][6] , \DataMem/Mem[1][7] ,
         \DataMem/Mem[1][8] , \DataMem/Mem[1][9] , \DataMem/Mem[1][10] ,
         \DataMem/Mem[1][11] , \DataMem/Mem[1][12] , \DataMem/Mem[1][13] ,
         \DataMem/Mem[1][14] , \DataMem/Mem[1][15] , \DataMem/Mem[1][16] ,
         \DataMem/Mem[1][17] , \DataMem/Mem[1][18] , \DataMem/Mem[1][19] ,
         \DataMem/Mem[1][20] , \DataMem/Mem[1][21] , \DataMem/Mem[1][22] ,
         \DataMem/Mem[1][23] , \DataMem/Mem[1][24] , \DataMem/Mem[1][25] ,
         \DataMem/Mem[1][26] , \DataMem/Mem[1][27] , \DataMem/Mem[1][28] ,
         \DataMem/Mem[1][29] , \DataMem/Mem[1][30] , \DataMem/Mem[1][31] ,
         \DataMem/Mem[2][0] , \DataMem/Mem[2][1] , \DataMem/Mem[2][2] ,
         \DataMem/Mem[2][3] , \DataMem/Mem[2][4] , \DataMem/Mem[2][5] ,
         \DataMem/Mem[2][6] , \DataMem/Mem[2][7] , \DataMem/Mem[2][8] ,
         \DataMem/Mem[2][9] , \DataMem/Mem[2][10] , \DataMem/Mem[2][11] ,
         \DataMem/Mem[2][12] , \DataMem/Mem[2][13] , \DataMem/Mem[2][14] ,
         \DataMem/Mem[2][15] , \DataMem/Mem[2][16] , \DataMem/Mem[2][17] ,
         \DataMem/Mem[2][18] , \DataMem/Mem[2][19] , \DataMem/Mem[2][20] ,
         \DataMem/Mem[2][21] , \DataMem/Mem[2][22] , \DataMem/Mem[2][23] ,
         \DataMem/Mem[2][24] , \DataMem/Mem[2][25] , \DataMem/Mem[2][26] ,
         \DataMem/Mem[2][27] , \DataMem/Mem[2][28] , \DataMem/Mem[2][29] ,
         \DataMem/Mem[2][30] , \DataMem/Mem[2][31] , \DataMem/Mem[3][0] ,
         \DataMem/Mem[3][1] , \DataMem/Mem[3][2] , \DataMem/Mem[3][3] ,
         \DataMem/Mem[3][4] , \DataMem/Mem[3][5] , \DataMem/Mem[3][6] ,
         \DataMem/Mem[3][7] , \DataMem/Mem[3][8] , \DataMem/Mem[3][9] ,
         \DataMem/Mem[3][10] , \DataMem/Mem[3][11] , \DataMem/Mem[3][12] ,
         \DataMem/Mem[3][13] , \DataMem/Mem[3][14] , \DataMem/Mem[3][15] ,
         \DataMem/Mem[3][16] , \DataMem/Mem[3][17] , \DataMem/Mem[3][18] ,
         \DataMem/Mem[3][19] , \DataMem/Mem[3][20] , \DataMem/Mem[3][21] ,
         \DataMem/Mem[3][22] , \DataMem/Mem[3][23] , \DataMem/Mem[3][24] ,
         \DataMem/Mem[3][25] , \DataMem/Mem[3][26] , \DataMem/Mem[3][27] ,
         \DataMem/Mem[3][28] , \DataMem/Mem[3][29] , \DataMem/Mem[3][30] ,
         \DataMem/Mem[3][31] , \DataMem/Mem[4][0] , \DataMem/Mem[4][1] ,
         \DataMem/Mem[4][2] , \DataMem/Mem[4][3] , \DataMem/Mem[4][4] ,
         \DataMem/Mem[4][5] , \DataMem/Mem[4][6] , \DataMem/Mem[4][7] ,
         \DataMem/Mem[4][8] , \DataMem/Mem[4][9] , \DataMem/Mem[4][10] ,
         \DataMem/Mem[4][11] , \DataMem/Mem[4][12] , \DataMem/Mem[4][13] ,
         \DataMem/Mem[4][14] , \DataMem/Mem[4][15] , \DataMem/Mem[4][16] ,
         \DataMem/Mem[4][17] , \DataMem/Mem[4][18] , \DataMem/Mem[4][19] ,
         \DataMem/Mem[4][20] , \DataMem/Mem[4][21] , \DataMem/Mem[4][22] ,
         \DataMem/Mem[4][23] , \DataMem/Mem[4][24] , \DataMem/Mem[4][25] ,
         \DataMem/Mem[4][26] , \DataMem/Mem[4][27] , \DataMem/Mem[4][28] ,
         \DataMem/Mem[4][29] , \DataMem/Mem[4][30] , \DataMem/Mem[4][31] ,
         \DataMem/Mem[5][0] , \DataMem/Mem[5][1] , \DataMem/Mem[5][2] ,
         \DataMem/Mem[5][3] , \DataMem/Mem[5][4] , \DataMem/Mem[5][5] ,
         \DataMem/Mem[5][6] , \DataMem/Mem[5][7] , \DataMem/Mem[5][8] ,
         \DataMem/Mem[5][9] , \DataMem/Mem[5][10] , \DataMem/Mem[5][11] ,
         \DataMem/Mem[5][12] , \DataMem/Mem[5][13] , \DataMem/Mem[5][14] ,
         \DataMem/Mem[5][15] , \DataMem/Mem[5][16] , \DataMem/Mem[5][17] ,
         \DataMem/Mem[5][18] , \DataMem/Mem[5][19] , \DataMem/Mem[5][20] ,
         \DataMem/Mem[5][21] , \DataMem/Mem[5][22] , \DataMem/Mem[5][23] ,
         \DataMem/Mem[5][24] , \DataMem/Mem[5][25] , \DataMem/Mem[5][26] ,
         \DataMem/Mem[5][27] , \DataMem/Mem[5][28] , \DataMem/Mem[5][29] ,
         \DataMem/Mem[5][30] , \DataMem/Mem[5][31] , \DataMem/Mem[6][0] ,
         \DataMem/Mem[6][1] , \DataMem/Mem[6][2] , \DataMem/Mem[6][3] ,
         \DataMem/Mem[6][4] , \DataMem/Mem[6][5] , \DataMem/Mem[6][6] ,
         \DataMem/Mem[6][7] , \DataMem/Mem[6][8] , \DataMem/Mem[6][9] ,
         \DataMem/Mem[6][10] , \DataMem/Mem[6][11] , \DataMem/Mem[6][12] ,
         \DataMem/Mem[6][13] , \DataMem/Mem[6][14] , \DataMem/Mem[6][15] ,
         \DataMem/Mem[6][16] , \DataMem/Mem[6][17] , \DataMem/Mem[6][18] ,
         \DataMem/Mem[6][19] , \DataMem/Mem[6][20] , \DataMem/Mem[6][21] ,
         \DataMem/Mem[6][22] , \DataMem/Mem[6][23] , \DataMem/Mem[6][24] ,
         \DataMem/Mem[6][25] , \DataMem/Mem[6][26] , \DataMem/Mem[6][27] ,
         \DataMem/Mem[6][28] , \DataMem/Mem[6][29] , \DataMem/Mem[6][30] ,
         \DataMem/Mem[6][31] , \DataMem/Mem[7][0] , \DataMem/Mem[7][1] ,
         \DataMem/Mem[7][2] , \DataMem/Mem[7][3] , \DataMem/Mem[7][4] ,
         \DataMem/Mem[7][5] , \DataMem/Mem[7][6] , \DataMem/Mem[7][7] ,
         \DataMem/Mem[7][8] , \DataMem/Mem[7][9] , \DataMem/Mem[7][10] ,
         \DataMem/Mem[7][11] , \DataMem/Mem[7][12] , \DataMem/Mem[7][13] ,
         \DataMem/Mem[7][14] , \DataMem/Mem[7][15] , \DataMem/Mem[7][16] ,
         \DataMem/Mem[7][17] , \DataMem/Mem[7][18] , \DataMem/Mem[7][19] ,
         \DataMem/Mem[7][20] , \DataMem/Mem[7][21] , \DataMem/Mem[7][22] ,
         \DataMem/Mem[7][23] , \DataMem/Mem[7][24] , \DataMem/Mem[7][25] ,
         \DataMem/Mem[7][26] , \DataMem/Mem[7][27] , \DataMem/Mem[7][28] ,
         \DataMem/Mem[7][29] , \DataMem/Mem[7][30] , \DataMem/Mem[7][31] ,
         \DataMem/N31 , \DataMem/N30 , \DataMem/N29 , \DataMem/N28 ,
         \DataMem/N27 , \DataMem/N26 , \DataMem/N25 , \DataMem/N24 ,
         \DataMem/N23 , \DataMem/N22 , \DataMem/N21 , \DataMem/N20 ,
         \DataMem/N19 , \DataMem/N18 , \DataMem/N17 , \DataMem/N16 ,
         \DataMem/N15 , \DataMem/N14 , \DataMem/N13 , \DataMem/N12 ,
         \DataMem/N11 , \DataMem/N10 , \DataMem/N9 , \DataMem/N8 ,
         \DataMem/N7 , \DataMem/N6 , \DataMem/N5 , \DataMem/N4 , \DataMem/N3 ,
         \DataMem/N2 , \DataMem/N1 , \DataMem/N0 , n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n4376, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7709, n7710, n7711, net175543, n12649,
         n12766, n13055, n13058, n13061, n13064, n13067, n13070, n13073,
         n13076, n13079, n13082, n13085, n13088, n13091, n13094, n13097,
         n13100, n13103, n13106, n13109, n13112, n13115, n13118, n13121,
         n13124, n13127, n13130, n13133, n13136, n13139, n13142, n13145,
         n13148, n13151, n13154, n13157, n13160, n13163, n13166, n13169,
         n13172, n13175, n13178, n13181, n13184, n13187, n13190, n13193,
         n13196, n13199, n13202, n13205, n13208, n13211, n13214, n13217,
         n13220, n13223, n13226, n13229, n13232, n13235, n13238, n13241,
         n13244, n13247, n13250, n13253, n13256, n13259, n13262, n13265,
         n13268, n13281, n13782, n13783, n13784, n13785, n13786, n13787,
         n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
         n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
         n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
         n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
         n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
         n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
         n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
         n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
         n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875,
         n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
         n13884, n13885, n13886, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13936, n13937, n13938,
         n13939, n13940, n13942, n13944, n13945, n13946, n13947, n13948,
         n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956,
         n13957, n13958, n13959, n13960, n13962, n13963, n13964, n13965,
         n13966, n13967, n13969, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14040, n14041, n14042, n14043, n14044,
         n14045, n14046, n14047, n14048, n14049, n14051, n14053, n14058,
         n14059, n14061, n14064, n14065, n14066, n14067, n14068, n14069,
         n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
         n14078, n14082, n14083, n14084, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14113, n14116, n14117, n14119, n14120, n14121, n14122, n14123,
         n14125, n14126, n14127, n14129, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14172, n14173, n14174, n14176, n14177, n14178,
         n14179, n14180, n14181, n14183, n14184, n14185, n14186, n14187,
         n14188, n14189, n14190, n14200, n14201, n14202, n14203, n14204,
         n14205, n14206, n14207, n14208, n14210, n14212, n14213, n14214,
         n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222,
         n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230,
         n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238,
         n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246,
         n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254,
         n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262,
         n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270,
         n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278,
         n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286,
         n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294,
         n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302,
         n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310,
         n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318,
         n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326,
         n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334,
         n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342,
         n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350,
         n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358,
         n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366,
         n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374,
         n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382,
         n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390,
         n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398,
         n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406,
         n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414,
         n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422,
         n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430,
         n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438,
         n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446,
         n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454,
         n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462,
         n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470,
         n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478,
         n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486,
         n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494,
         n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502,
         n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510,
         n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518,
         n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526,
         n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534,
         n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542,
         n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550,
         n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558,
         n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566,
         n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574,
         n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582,
         n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590,
         n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598,
         n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606,
         n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614,
         n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622,
         n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630,
         n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638,
         n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646,
         n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654,
         n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662,
         n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670,
         n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678,
         n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686,
         n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694,
         n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702,
         n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710,
         n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718,
         n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726,
         n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734,
         n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742,
         n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750,
         n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758,
         n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766,
         n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774,
         n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782,
         n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790,
         n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798,
         n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806,
         n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814,
         n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822,
         n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830,
         n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838,
         n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846,
         n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854,
         n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862,
         n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870,
         n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878,
         n14879, n14880, n14881, n14882, n14883, n14885, n14887, n14889,
         n14891, n14893, n14895, n14897, n14899, n14901, n14903, n14905,
         n14907, n14909, n14911, n14913, n14915, n14917, n14919, n14921,
         n14923, n14925, n14927, n14929, n14931, n14933, n14935, n14937,
         n14939, n14941, n14943, n14945, n14947, n14948, n14949, n14950,
         n14951, n14952, n14954, n14955, n14956, n14957, n14958, n14959,
         n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967,
         n14968, n14970, n14971, n14972, n14974, n14975, n14976, n14977,
         n14978, n14979, n14981, n14982, n14988, n14993, n14995, n15001,
         n15007, n15009, n15010, n15011, n15013, n15014, n15015, n15017,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15029, n15030, n15032, n15033, n15034, n15035, n15037, n15039,
         n15040, n15041, n15042, n15043, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15062, n15064, n15066, n15068, n15070, n15072,
         n15074, n15076, n15078, n15080, n15082, n15084, n15086, n15088,
         n15090, n15092, n15094, n15096, n15098, n15100, n15102, n15104,
         n15106, n15108, n15110, n15112, n15114, n15116, n15118, n15120,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15133, n15134, n15137, n15138, n15142, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15180, n15181,
         n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189,
         n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198,
         n15199, n15201, n15202, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15233, n15234,
         n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
         n15243, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
         n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15260,
         n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268,
         n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276,
         n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285,
         n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15294,
         n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302,
         n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15311,
         n15312, n15313, n15314, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15345, n15346,
         n15348, n15352, n15353, n15354, n15355, n15356, n15357, n15358,
         n15359, n15360, n15362, n15363, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15381, n15382, n15383, n15384, n15385, n15386,
         n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15395,
         n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403,
         n15404, n15405, n15406, n15407, n15408, n15410, n15411, n15412,
         n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420,
         n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428,
         n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436,
         n15437, n15438, n15439, n15440, n15441, n15442, n15444, n15445,
         n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453,
         n15454, n15455, n15456, n15458, n15459, n15460, n15461, n15462,
         n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470,
         n15471, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
         n15480, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514,
         n15515, n15516, n15517, n15518, n15519, n15521, n15522, n15523,
         n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531,
         n15532, n15533, n15534, n15535, n15537, n15538, n15539, n15540,
         n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548,
         n15549, n15550, n15552, n15553, n15554, n15555, n15556, n15557,
         n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15566,
         n15567, n15568, n15569, n15570, n15571, n15573, n15574, n15575,
         n15576, n15577, n15578, n15579, n15581, n15582, n15583, n15584,
         n15586, n15588, n15590, n15591, n15592, n15593, n15594, n15595,
         n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603,
         n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611,
         n15612, n15621, n15622, n15623, n15624, n15625, n15626, n15627,
         n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635,
         n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643,
         n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651,
         n15652, n15653, n15686, n15687, n15688, n15689, n15690, n15691,
         n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699,
         n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707,
         n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715,
         n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723,
         n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731,
         n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739,
         n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747,
         n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755,
         n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763,
         n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771,
         n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779,
         n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787,
         n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795,
         n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803,
         n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811,
         n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819,
         n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827,
         n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835,
         n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843,
         n15844, n15845, n15846, n15847, n15848, n15849, n15866, n15867,
         n15868, n15869, n15886, n15887, n15888, n15889, n15890, n15891,
         n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899,
         n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908,
         n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916,
         n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924,
         n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932,
         n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940,
         n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948,
         n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956,
         n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964,
         n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972,
         n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980,
         n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988,
         n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996,
         n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004,
         n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012,
         n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020,
         n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028,
         n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036,
         n16037, n16038, n16039, n16040, n16041, n16042, n16043, n16044,
         n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052,
         n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060,
         n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068,
         n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076,
         n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084,
         n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092,
         n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100,
         n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108,
         n16109, n16110, n16111, n16112, n16113, n16114, n16115, n16116,
         n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124,
         n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132,
         n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140,
         n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148,
         n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156,
         n16157, n16158, n16159, n16160, n16161, n16162, n16163, n16164,
         n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172,
         n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180,
         n16181, n16182, n16183, n16184, n16185, n16186, n16187, n16188,
         n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196,
         n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204,
         n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212,
         n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220,
         n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228,
         n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236,
         n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244,
         n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252,
         n16253, n16254, n16255, n16256, n16257, n16258, n16259, n16260,
         n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268,
         n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276,
         n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284,
         n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292,
         n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300,
         n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308,
         n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316,
         n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324,
         n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332,
         n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340,
         n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348,
         n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356,
         n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364,
         n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372,
         n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380,
         n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388,
         n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396,
         n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404,
         n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412,
         n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420,
         n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428,
         n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436,
         n16437, n16438, n16439, n16440, n16441, n16442, n16443, n16444,
         n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452,
         n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460,
         n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468,
         n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476,
         n16477, n16478, n16479, n16480, n16481, n16482, n16483, n16484,
         n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492,
         n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500,
         n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508,
         n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516,
         n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524,
         n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532,
         n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540,
         n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548,
         n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556,
         n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16565,
         n16568, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16603, n16605,
         n16606, n16607, n16608, n16609, n16611, n16612, n16614, n16615,
         n16616, n16617, n16618, n16619, n16620, n16624, n16626, n16629,
         n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637,
         n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645,
         n16646, n16647, n16648, n16649, n16650, n16651, n16652, n16653,
         n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661,
         n16662, n16663, n16664, n16666, n16667, n16668, n16669, n16670,
         n16671, n16672, n16676, n16677, n16678, n16679, n16680, n16681,
         n16683, n16684, n16685, n16686, n16687, n16689, n16690, n16691,
         n16693, n16696, n16699, n16701, n16704, n16710, n16711, n16712,
         n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720,
         n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728,
         n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736,
         n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744,
         n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752,
         n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760,
         n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768,
         n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776,
         n16777, n16778, n16779, n16780, n16784, n16785, n16786, n16789,
         n16790, n16791, n16792, n16793, n16795, n16796, n16806, n16807,
         n16808, n16809, n16811, n16812, n16813, n16814, n16815, n16816,
         n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824,
         n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832,
         n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840,
         n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848,
         n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856,
         n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864,
         n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872,
         n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880,
         n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888,
         n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896,
         n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904,
         n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912,
         n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920,
         n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928,
         n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936,
         n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944,
         n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952,
         n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960,
         n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968,
         n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976,
         n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984,
         n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992,
         n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000,
         n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008,
         n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016,
         n16613, n16682, n16688, n16805, n15000, n16783, n16782, n15005,
         \pipeline/stageF/PC_plus4/add_26/n1 ,
         \pipeline/stageF/PC_plus4/add_26/carry[4] ,
         \pipeline/stageF/PC_plus4/add_26/carry[5] ,
         \pipeline/stageF/PC_plus4/add_26/carry[6] ,
         \pipeline/stageF/PC_plus4/add_26/carry[7] ,
         \pipeline/stageF/PC_plus4/add_26/carry[8] ,
         \pipeline/stageF/PC_plus4/add_26/carry[9] ,
         \pipeline/stageF/PC_plus4/add_26/carry[10] ,
         \pipeline/stageF/PC_plus4/add_26/carry[11] ,
         \pipeline/stageF/PC_plus4/add_26/carry[12] ,
         \pipeline/stageF/PC_plus4/add_26/carry[13] ,
         \pipeline/stageF/PC_plus4/add_26/carry[14] ,
         \pipeline/stageF/PC_plus4/add_26/carry[15] ,
         \pipeline/stageF/PC_plus4/add_26/carry[16] ,
         \pipeline/stageF/PC_plus4/add_26/carry[17] ,
         \pipeline/stageF/PC_plus4/add_26/carry[18] ,
         \pipeline/stageF/PC_plus4/add_26/carry[19] ,
         \pipeline/stageF/PC_plus4/add_26/carry[20] ,
         \pipeline/stageF/PC_plus4/add_26/carry[21] ,
         \pipeline/stageF/PC_plus4/add_26/carry[22] ,
         \pipeline/stageF/PC_plus4/add_26/carry[23] ,
         \pipeline/stageF/PC_plus4/add_26/carry[24] ,
         \pipeline/stageF/PC_plus4/add_26/carry[25] ,
         \pipeline/stageF/PC_plus4/add_26/carry[26] ,
         \pipeline/stageF/PC_plus4/add_26/carry[27] ,
         \pipeline/stageF/PC_plus4/add_26/carry[28] ,
         \pipeline/stageF/PC_plus4/add_26/carry[29] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n170 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n169 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n167 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n166 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n165 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n164 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n163 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n162 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n161 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n160 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n158 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n157 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n156 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n155 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n154 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n153 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n152 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n151 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n150 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n149 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n148 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n145 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n144 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n143 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n140 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n139 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n136 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n135 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n134 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n133 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n132 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n127 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n124 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n121 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n118 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n117 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n116 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n115 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n114 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n113 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n112 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n111 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n110 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n109 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n108 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n107 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n106 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n105 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n103 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n102 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n101 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n100 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n99 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n98 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n94 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n93 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n92 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n91 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n90 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n89 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n88 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n87 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n86 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n85 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n84 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n83 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n82 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n81 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n80 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n79 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n78 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n77 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n76 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n75 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n74 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n73 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n72 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n71 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n70 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n69 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n68 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n67 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n66 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n64 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n63 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n62 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n61 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n60 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n59 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n58 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n56 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n54 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n53 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n52 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n51 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n50 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n48 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n46 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n45 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n44 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n43 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n42 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n41 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n40 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n39 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n38 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n37 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n36 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n35 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n34 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n33 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n32 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n31 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n30 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n29 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n28 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n27 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n26 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n25 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n24 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n23 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n22 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n21 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n20 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n19 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n18 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n17 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n16 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n15 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n14 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n13 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n12 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n11 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n10 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n9 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n8 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n7 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n6 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n5 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n4 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n2 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/n1 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[1] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[3] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C48/A[16] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n172 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n171 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n170 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n169 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n168 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n167 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n165 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n163 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n162 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n161 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n160 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n158 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n156 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n154 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n153 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n152 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n149 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n146 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n144 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n143 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n142 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n140 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n139 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n138 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n136 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n135 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n134 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n133 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n131 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n130 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n129 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n128 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n127 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n126 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n122 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n121 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n120 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n118 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n117 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n116 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n114 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n113 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n112 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n111 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n109 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n108 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n107 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n106 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n104 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n103 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n102 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n101 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n99 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n98 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n97 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n96 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n95 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n94 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n92 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n91 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n90 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n89 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n88 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n87 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n85 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n84 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n83 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n82 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n81 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n80 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n79 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n77 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n76 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n75 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n74 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n73 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n72 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n71 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n70 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n69 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n68 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n67 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n66 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n64 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n63 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n62 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n61 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n60 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n58 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n57 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n56 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n55 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n54 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n53 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n52 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n50 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n49 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n48 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n47 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n46 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n45 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n44 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n42 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n41 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n40 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n39 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n38 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n37 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n36 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n35 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n33 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n32 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n31 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n30 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n29 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n28 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n27 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n26 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n25 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n23 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n21 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n20 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n19 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n18 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n17 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n16 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n15 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n14 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n13 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n12 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n11 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n10 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n9 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n8 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n7 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n6 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n5 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n4 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n3 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C86/n1 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][0] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][1] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][2] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][3] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][4] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][5] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][6] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][7] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][8] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][9] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][10] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][11] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][12] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][13] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][14] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][15] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][16] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][17] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][18] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][19] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][20] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][21] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][22] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][23] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][24] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][25] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][26] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][27] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][28] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][29] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][30] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][31] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][0] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][1] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][2] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][3] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][4] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][5] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][6] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][7] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][8] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][9] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][10] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][11] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][12] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][13] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][14] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][15] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][16] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][17] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][18] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][19] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][20] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][21] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][22] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][23] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][24] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][25] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][26] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][27] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][28] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][29] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][30] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][31] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][0] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][1] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][2] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][3] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][4] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][5] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][6] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][7] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][8] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][9] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][10] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][11] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][12] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][13] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][14] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][15] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][16] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][17] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][18] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][19] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][20] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][21] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][22] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][23] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][24] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][25] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][26] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][27] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][28] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][29] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][30] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][31] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][0] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][1] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][2] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][3] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][5] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][6] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][7] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][8] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][9] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][10] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][11] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][12] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][13] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][14] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][15] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][16] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][17] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][18] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][19] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][20] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][21] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][22] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][23] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][24] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][25] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][26] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][27] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][28] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][29] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][30] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][31] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][0] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][1] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][2] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][3] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][4] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][5] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][6] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][7] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][8] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][9] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][10] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][11] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][12] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][13] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][14] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][15] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][16] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][17] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][18] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][19] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][20] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][21] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][22] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][23] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][24] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][25] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][26] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][27] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][28] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][29] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][30] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][31] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][0] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][1] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][2] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][3] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][4] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][5] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][6] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][7] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][8] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][9] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][10] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][11] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][12] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][13] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][14] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][15] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][16] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][17] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][18] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][19] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][20] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][21] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][22] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][23] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][24] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][25] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][26] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][27] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][28] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][29] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][30] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][31] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][0] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][1] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][2] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][3] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][4] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][5] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][6] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][7] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][8] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][9] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][10] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][11] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][12] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][13] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][14] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][15] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][16] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][17] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][18] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][19] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][20] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][21] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][22] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][23] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][24] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][25] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][26] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][27] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][28] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][29] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][30] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][31] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][0] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][1] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][2] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][3] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][4] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][5] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][6] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][7] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][8] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][9] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][10] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][11] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][12] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][13] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][14] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][15] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][16] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][17] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][18] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][19] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][20] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][21] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][22] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][23] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][24] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][25] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][26] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][27] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][28] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][29] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][30] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][31] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n167 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n161 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n160 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n159 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n158 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n157 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n156 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n155 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n153 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n151 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n148 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n147 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n146 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n145 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n144 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n143 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n142 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n141 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n139 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n138 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n137 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n132 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n131 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n128 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n127 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n126 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n125 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n124 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n123 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n122 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n121 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n120 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n117 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n114 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n108 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n105 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n104 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n103 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n102 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n101 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n100 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n99 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n98 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n97 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n96 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n95 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n94 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n93 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n92 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n91 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n90 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n89 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n88 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n87 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n83 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n82 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n81 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n80 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n79 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n78 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n77 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n76 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n75 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n74 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n73 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n72 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n71 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n70 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n69 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n68 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n67 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n66 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n65 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n63 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n62 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n61 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n60 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n59 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n58 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n57 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n55 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n53 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n51 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n50 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n49 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n48 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n46 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n44 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n43 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n42 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n41 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n40 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n39 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n38 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n37 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n36 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n35 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n34 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n33 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n32 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n31 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n30 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n29 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n28 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n27 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n26 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n25 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n24 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n23 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n22 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n21 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n20 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n19 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n18 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n17 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n16 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n15 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n14 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n13 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n12 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n11 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n10 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n9 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n8 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n7 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n6 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n5 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n4 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n3 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C50/n2 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/n10 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/n9 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/n8 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/n7 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/n6 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/n5 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/n4 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/n3 ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][0] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][1] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][2] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][3] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][4] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][5] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][6] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][7] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][8] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][9] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][10] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][11] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][12] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][13] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][14] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][15] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][16] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][17] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][18] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][19] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][20] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][21] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][22] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][23] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][24] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][25] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][26] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][27] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][28] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][29] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][30] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][31] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][0] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][1] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][2] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][3] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][4] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][5] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][6] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][7] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][8] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][9] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][10] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][11] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][12] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][13] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][14] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][15] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][16] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][17] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][18] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][19] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][20] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][21] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][22] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][23] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][24] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][25] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][26] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][27] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][28] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][29] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][30] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][31] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][0] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][1] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][2] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][3] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][4] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][5] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][6] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][7] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][8] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][9] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][10] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][11] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][12] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][13] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][14] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][15] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][16] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][17] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][18] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][19] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][20] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][21] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][22] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][23] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][24] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][25] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][26] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][27] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][28] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][29] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][30] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][31] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][0] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][1] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][2] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][3] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][4] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][5] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][6] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][7] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][8] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][9] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][10] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][11] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][12] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][13] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][14] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][15] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][16] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][17] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][18] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][19] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][20] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][21] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][22] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][23] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][24] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][25] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][26] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][27] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][28] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][29] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][30] ,
         \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][31] ,
         \pipeline/stageD/evaluate_jump_target/add_29/n214 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n213 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n209 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n208 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n207 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n203 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n202 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n201 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n197 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n196 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n195 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n194 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n191 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n190 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n189 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n188 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n185 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n184 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n183 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n182 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n181 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n180 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n178 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n177 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n175 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n174 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n172 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n171 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n170 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n169 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n168 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n165 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n163 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n160 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n159 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n157 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n150 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n149 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n145 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n144 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n141 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n139 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n138 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n135 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n134 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n133 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n132 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n129 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n128 ,
         \pipeline/stageD/evaluate_jump_target/add_29/n126 , n17018, n17019,
         n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027,
         n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035,
         n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043,
         n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051,
         n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059,
         n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067,
         n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075,
         n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083,
         n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091,
         n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099,
         n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107,
         n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115,
         n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123,
         n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131,
         n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139,
         n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147,
         n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155,
         n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163,
         n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171,
         n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179,
         n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187,
         n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195,
         n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203,
         n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211,
         n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219,
         n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227,
         n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235,
         n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243,
         n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251,
         n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259,
         n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267,
         n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275,
         n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283,
         n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291,
         n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299,
         n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307,
         n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315,
         n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323,
         n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331,
         n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339,
         n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347,
         n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355,
         n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363,
         n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371,
         n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379,
         n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387,
         n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395,
         n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403,
         n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411,
         n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419,
         n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427,
         n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435,
         n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443,
         n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451,
         n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459,
         n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467,
         n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475,
         n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483,
         n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491,
         n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499,
         n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507,
         n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515,
         n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523,
         n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531,
         n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539,
         n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547,
         n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555,
         n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563,
         n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571,
         n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579,
         n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587,
         n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595,
         n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603,
         n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611,
         n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619,
         n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627,
         n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635,
         n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643,
         n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651,
         n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659,
         n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667,
         n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675,
         n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683,
         n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691,
         n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699,
         n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707,
         n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715,
         n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723,
         n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731,
         n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739,
         n17740, n17741, n17742, n17743, n17744;
  wire   [31:0] InstrFetched;
  wire   [31:0] addr_to_dataRam;
  wire   [31:0] \pipeline/immediate_to_exe ;
  wire   [4:0] \pipeline/Reg2_Addr_to_exe ;
  wire   [4:0] \pipeline/Reg1_Addr_to_exe ;
  wire   [8:0] \pipeline/EXE_controls_in_EXEcute ;
  wire   [31:0] \pipeline/stageD/offset_to_jump_temp ;
  wire   [31:0] \pipeline/stageD/offset_jump_sign_ext ;
  wire   [31:0] \pipeline/stageE/input1_to_ALU ;
  tri   [31:0] addr_to_iram;
  tri   [31:0] data_from_dram;
  tri   \pipeline/stageF/PC_plus4/N8 ;
  tri   \pipeline/stageF/PC_plus4/N7 ;
  tri   [31:0] \pipeline/stageD/target_Jump_temp ;
  assign n13281 = Rst;

  DLH_X1 \DataMem/Mem_reg[7][31]  ( .G(n13079), .D(\DataMem/N2159 ), .Q(
        \DataMem/Mem[7][31] ) );
  DLL_X1 \DataMem/Dataout_reg[31]  ( .D(\DataMem/N2254 ), .GN(n17098), .Q(
        \DataMem/N2256 ) );
  DFF_X1 \pipeline/MEMWB_Stage/Data_to_RF_reg[31]  ( .D(
        \pipeline/MEMWB_Stage/N42 ), .CK(Clk), .Q(
        \pipeline/data_to_RF_from_WB[31] ), .QN(n17425) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[1][31]  ( .G(n13172), .D(n13268), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[1][31] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg1_out_IDEX_reg[31]  ( .D(
        \pipeline/IDEX_Stage/N133 ), .CK(Clk), .Q(n13966) );
  DFF_X1 \pipeline/MEMWB_Stage/Data_to_RF_reg[0]  ( .D(
        \pipeline/MEMWB_Stage/N11 ), .CK(Clk), .Q(
        \pipeline/data_to_RF_from_WB[0] ), .QN(n17396) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[1][0]  ( .G(n17706), .D(n13175), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[1][0] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg1_out_IDEX_reg[0]  ( .D(
        \pipeline/IDEX_Stage/N102 ), .CK(Clk), .Q(n13965) );
  DFF_X1 \pipeline/MEMWB_Stage/Data_to_RF_reg[8]  ( .D(
        \pipeline/MEMWB_Stage/N19 ), .CK(Clk), .Q(
        \pipeline/data_to_RF_from_WB[8] ), .QN(n17394) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[1][8]  ( .G(n17706), .D(n13199), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[1][8] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg1_out_IDEX_reg[8]  ( .D(
        \pipeline/IDEX_Stage/N110 ), .CK(Clk), .Q(n13964) );
  DFF_X1 \pipeline/MEMWB_Stage/Data_to_RF_reg[24]  ( .D(
        \pipeline/MEMWB_Stage/N35 ), .CK(Clk), .Q(
        \pipeline/data_to_RF_from_WB[24] ), .QN(n17324) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[1][24]  ( .G(n13172), .D(n13247), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[1][24] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg1_out_IDEX_reg[24]  ( .D(
        \pipeline/IDEX_Stage/N126 ), .CK(Clk), .Q(n13963) );
  DFF_X1 \pipeline/MEMWB_Stage/Data_to_RF_reg[28]  ( .D(
        \pipeline/MEMWB_Stage/N39 ), .CK(Clk), .Q(
        \pipeline/data_to_RF_from_WB[28] ), .QN(n17312) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[1][28]  ( .G(n13172), .D(n13259), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[1][28] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg1_out_IDEX_reg[28]  ( .D(
        \pipeline/IDEX_Stage/N130 ), .CK(Clk), .Q(n13962) );
  DFF_X1 \pipeline/IFID_stage/Instr_out_IFID_reg[14]  ( .D(n3992), .CK(Clk), 
        .Q(\pipeline/stageD/offset_to_jump_temp [14]), .QN(n17445) );
  DFF_X1 \pipeline/IDEX_Stage/Immediate_out_IDEX_reg[14]  ( .D(
        \pipeline/IDEX_Stage/N180 ), .CK(Clk), .Q(
        \pipeline/immediate_to_exe [14]) );
  DFF_X1 \pipeline/MEMWB_Stage/Data_to_RF_reg[14]  ( .D(
        \pipeline/MEMWB_Stage/N25 ), .CK(Clk), .Q(
        \pipeline/data_to_RF_from_WB[14] ), .QN(n17309) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[1][14]  ( .G(n13172), .D(n13217), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[1][14] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg1_out_IDEX_reg[14]  ( .D(
        \pipeline/IDEX_Stage/N116 ), .CK(Clk), .Q(n13960) );
  DFF_X1 \pipeline/MEMWB_Stage/Data_to_RF_reg[15]  ( .D(
        \pipeline/MEMWB_Stage/N26 ), .CK(Clk), .Q(
        \pipeline/data_to_RF_from_WB[15] ), .QN(n17364) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[1][15]  ( .G(n17706), .D(n13220), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[1][15] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg1_out_IDEX_reg[15]  ( .D(
        \pipeline/IDEX_Stage/N117 ), .CK(Clk), .Q(n13959) );
  DFF_X1 \pipeline/MEMWB_Stage/Data_to_RF_reg[13]  ( .D(
        \pipeline/MEMWB_Stage/N24 ), .CK(Clk), .Q(
        \pipeline/data_to_RF_from_WB[13] ), .QN(n17344) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[1][13]  ( .G(n13172), .D(n13214), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[1][13] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg1_out_IDEX_reg[13]  ( .D(
        \pipeline/IDEX_Stage/N115 ), .CK(Clk), .Q(n13958) );
  DFF_X1 \pipeline/MEMWB_Stage/Data_to_RF_reg[30]  ( .D(
        \pipeline/MEMWB_Stage/N41 ), .CK(Clk), .Q(
        \pipeline/data_to_RF_from_WB[30] ), .QN(n17362) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[1][30]  ( .G(n17706), .D(n13265), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[1][30] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg1_out_IDEX_reg[30]  ( .D(
        \pipeline/IDEX_Stage/N132 ), .CK(Clk), .Q(n13957) );
  DFF_X1 \pipeline/MEMWB_Stage/Data_to_RF_reg[29]  ( .D(
        \pipeline/MEMWB_Stage/N40 ), .CK(Clk), .Q(
        \pipeline/data_to_RF_from_WB[29] ), .QN(n17365) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[1][29]  ( .G(n17706), .D(n13262), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[1][29] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg1_out_IDEX_reg[29]  ( .D(
        \pipeline/IDEX_Stage/N131 ), .CK(Clk), .Q(n13956) );
  DFF_X1 \pipeline/MEMWB_Stage/Data_to_RF_reg[27]  ( .D(
        \pipeline/MEMWB_Stage/N38 ), .CK(Clk), .Q(
        \pipeline/data_to_RF_from_WB[27] ), .QN(n17325) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[1][27]  ( .G(n13172), .D(n13256), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[1][27] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg1_out_IDEX_reg[27]  ( .D(
        \pipeline/IDEX_Stage/N129 ), .CK(Clk), .Q(n13955) );
  DFF_X1 \pipeline/MEMWB_Stage/Data_to_RF_reg[26]  ( .D(
        \pipeline/MEMWB_Stage/N37 ), .CK(Clk), .Q(
        \pipeline/data_to_RF_from_WB[26] ), .QN(n17424) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[1][26]  ( .G(n13172), .D(n13253), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[1][26] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg1_out_IDEX_reg[26]  ( .D(
        \pipeline/IDEX_Stage/N128 ), .CK(Clk), .Q(n13954) );
  DFF_X1 \pipeline/MEMWB_Stage/Data_to_RF_reg[25]  ( .D(
        \pipeline/MEMWB_Stage/N36 ), .CK(Clk), .Q(
        \pipeline/data_to_RF_from_WB[25] ), .QN(n17427) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[1][25]  ( .G(n17706), .D(n13250), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[1][25] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg1_out_IDEX_reg[25]  ( .D(
        \pipeline/IDEX_Stage/N127 ), .CK(Clk), .Q(n13953) );
  DFF_X1 \pipeline/MEMWB_Stage/Data_to_RF_reg[23]  ( .D(
        \pipeline/MEMWB_Stage/N34 ), .CK(Clk), .Q(
        \pipeline/data_to_RF_from_WB[23] ), .QN(n17366) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[1][23]  ( .G(n17706), .D(n13244), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[1][23] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg1_out_IDEX_reg[23]  ( .D(
        \pipeline/IDEX_Stage/N125 ), .CK(Clk), .Q(n13952) );
  DFF_X1 \pipeline/MEMWB_Stage/Data_to_RF_reg[22]  ( .D(
        \pipeline/MEMWB_Stage/N33 ), .CK(Clk), .Q(
        \pipeline/data_to_RF_from_WB[22] ), .QN(n17311) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[1][22]  ( .G(n13172), .D(n13241), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[1][22] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg1_out_IDEX_reg[22]  ( .D(
        \pipeline/IDEX_Stage/N124 ), .CK(Clk), .Q(n13951) );
  DFF_X1 \pipeline/MEMWB_Stage/Data_to_RF_reg[21]  ( .D(
        \pipeline/MEMWB_Stage/N32 ), .CK(Clk), .Q(
        \pipeline/data_to_RF_from_WB[21] ), .QN(n17310) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[1][21]  ( .G(n13172), .D(n13238), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[1][21] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg1_out_IDEX_reg[21]  ( .D(
        \pipeline/IDEX_Stage/N123 ), .CK(Clk), .Q(n13950) );
  DFF_X1 \pipeline/MEMWB_Stage/Data_to_RF_reg[20]  ( .D(
        \pipeline/MEMWB_Stage/N31 ), .CK(Clk), .Q(
        \pipeline/data_to_RF_from_WB[20] ), .QN(n17322) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[1][20]  ( .G(n13172), .D(n13235), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[1][20] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg1_out_IDEX_reg[20]  ( .D(
        \pipeline/IDEX_Stage/N122 ), .CK(Clk), .Q(n13949) );
  DFF_X1 \pipeline/MEMWB_Stage/Data_to_RF_reg[19]  ( .D(
        \pipeline/MEMWB_Stage/N30 ), .CK(Clk), .Q(
        \pipeline/data_to_RF_from_WB[19] ), .QN(n17423) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[1][19]  ( .G(n17706), .D(n13232), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[1][19] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg1_out_IDEX_reg[19]  ( .D(
        \pipeline/IDEX_Stage/N121 ), .CK(Clk), .Q(n13948) );
  DFF_X1 \pipeline/MEMWB_Stage/Data_to_RF_reg[18]  ( .D(
        \pipeline/MEMWB_Stage/N29 ), .CK(Clk), .Q(
        \pipeline/data_to_RF_from_WB[18] ), .QN(n17363) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[1][18]  ( .G(n17706), .D(n13229), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[1][18] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg1_out_IDEX_reg[18]  ( .D(
        \pipeline/IDEX_Stage/N120 ), .CK(Clk), .Q(n13947) );
  DFF_X1 \pipeline/MEMWB_Stage/Data_to_RF_reg[17]  ( .D(
        \pipeline/MEMWB_Stage/N28 ), .CK(Clk), .Q(
        \pipeline/data_to_RF_from_WB[17] ), .QN(n17323) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[1][17]  ( .G(n13172), .D(n13226), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[1][17] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg1_out_IDEX_reg[17]  ( .D(
        \pipeline/IDEX_Stage/N119 ), .CK(Clk), .Q(n13946) );
  DFF_X1 \pipeline/MEMWB_Stage/Data_to_RF_reg[16]  ( .D(
        \pipeline/MEMWB_Stage/N27 ), .CK(Clk), .Q(
        \pipeline/data_to_RF_from_WB[16] ), .QN(n17426) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[1][16]  ( .G(n17706), .D(n13223), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[1][16] ) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_reg[16]  ( .D(n3991), .CK(Clk), .RN(
        n17704), .Q(n13945), .QN(n7711) );
  DFF_X1 \pipeline/IFID_stage/PC_out_IFID_reg[16]  ( .D(n3990), .CK(Clk), .Q(
        \pipeline/nextPC_IFID_DEC[16] ), .QN(n17461) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_reg[29]  ( .D(n3988), .CK(Clk), .RN(
        n17704), .Q(n13944), .QN(n7709) );
  DFF_X1 \pipeline/IFID_stage/Instr_out_IFID_reg[2]  ( .D(n3985), .CK(Clk), 
        .Q(\pipeline/stageD/offset_to_jump_temp [2]), .QN(n17404) );
  DFF_X1 \pipeline/IFID_stage/Instr_out_IFID_reg[3]  ( .D(n3984), .CK(Clk), 
        .Q(\pipeline/stageD/offset_to_jump_temp [3]), .QN(n17410) );
  DFF_X1 \pipeline/IFID_stage/Instr_out_IFID_reg[6]  ( .D(n3981), .CK(Clk), 
        .Q(\pipeline/stageD/offset_to_jump_temp [6]), .QN(n17361) );
  DFF_X1 \pipeline/IFID_stage/Instr_out_IFID_reg[7]  ( .D(n3980), .CK(Clk), 
        .Q(\pipeline/stageD/offset_to_jump_temp [7]), .QN(n17437) );
  DFF_X1 \pipeline/IFID_stage/Instr_out_IFID_reg[8]  ( .D(n3979), .CK(Clk), 
        .Q(\pipeline/stageD/offset_to_jump_temp [8]), .QN(n17428) );
  DFF_X1 \pipeline/IFID_stage/Instr_out_IFID_reg[9]  ( .D(n3978), .CK(Clk), 
        .Q(\pipeline/stageD/offset_to_jump_temp [9]), .QN(n17432) );
  DFF_X1 \pipeline/IFID_stage/Instr_out_IFID_reg[10]  ( .D(n3977), .CK(Clk), 
        .Q(\pipeline/stageD/offset_to_jump_temp [10]), .QN(n17440) );
  DFF_X1 \pipeline/IFID_stage/Instr_out_IFID_reg[11]  ( .D(n3976), .CK(Clk), 
        .Q(\pipeline/stageD/offset_to_jump_temp [11]), .QN(n17433) );
  DFF_X1 \pipeline/IFID_stage/Instr_out_IFID_reg[12]  ( .D(n3975), .CK(Clk), 
        .Q(\pipeline/stageD/offset_to_jump_temp [12]), .QN(n17444) );
  DFF_X1 \pipeline/IFID_stage/Instr_out_IFID_reg[13]  ( .D(n3974), .CK(Clk), 
        .Q(\pipeline/stageD/offset_to_jump_temp [13]), .QN(n17434) );
  DFF_X1 \pipeline/IFID_stage/Instr_out_IFID_reg[15]  ( .D(n3973), .CK(Clk), 
        .Q(\pipeline/stageD/offset_to_jump_temp [15]), .QN(n17431) );
  DFF_X1 \pipeline/IFID_stage/Instr_out_IFID_reg[16]  ( .D(n3972), .CK(Clk), 
        .Q(\pipeline/stageD/offset_jump_sign_ext [16]), .QN(n17316) );
  DFF_X1 \pipeline/IFID_stage/Instr_out_IFID_reg[17]  ( .D(n3971), .CK(Clk), 
        .Q(\pipeline/stageD/offset_jump_sign_ext [17]), .QN(n17329) );
  DFF_X1 \pipeline/IFID_stage/Instr_out_IFID_reg[18]  ( .D(n3970), .CK(Clk), 
        .Q(\pipeline/stageD/offset_jump_sign_ext [18]), .QN(n17408) );
  DFF_X1 \pipeline/IFID_stage/Instr_out_IFID_reg[19]  ( .D(n3969), .CK(Clk), 
        .Q(\pipeline/stageD/offset_jump_sign_ext [19]), .QN(n17349) );
  DFF_X1 \pipeline/IFID_stage/Instr_out_IFID_reg[20]  ( .D(n3968), .CK(Clk), 
        .Q(\pipeline/stageD/offset_jump_sign_ext [20]), .QN(n17407) );
  DFF_X1 \pipeline/IFID_stage/Instr_out_IFID_reg[26]  ( .D(n3962), .CK(Clk), 
        .Q(\pipeline/inst_IFID_DEC[26] ), .QN(n17409) );
  DFF_X1 \pipeline/IFID_stage/Instr_out_IFID_reg[28]  ( .D(n3960), .CK(Clk), 
        .Q(\pipeline/inst_IFID_DEC[28] ), .QN(n17348) );
  DFF_X1 \pipeline/IFID_stage/Instr_out_IFID_reg[30]  ( .D(n3958), .CK(Clk), 
        .Q(\pipeline/inst_IFID_DEC[30] ), .QN(n17347) );
  DLL_X1 \pipeline/cu_pipeline/ALU_OPCODE_reg[2]  ( .D(
        \pipeline/cu_pipeline/N103 ), .GN(n13281), .Q(
        \pipeline/EXE_controls_in_IDEX[3] ) );
  DLL_X1 \pipeline/cu_pipeline/ALU_OPCODE_reg[3]  ( .D(
        \pipeline/cu_pipeline/N104 ), .GN(n13281), .Q(
        \pipeline/EXE_controls_in_IDEX[4] ) );
  DLL_X1 \pipeline/cu_pipeline/ALU_OPCODE_reg[5]  ( .D(
        \pipeline/cu_pipeline/N106 ), .GN(n13281), .Q(
        \pipeline/EXE_controls_in_IDEX[6] ) );
  DLL_X1 \pipeline/cu_pipeline/ALU_OPCODE_reg[0]  ( .D(
        \pipeline/cu_pipeline/N101 ), .GN(n13281), .Q(
        \pipeline/EXE_controls_in_IDEX[1] ) );
  DLH_X1 \pipeline/cu_pipeline/Reg_dst_reg  ( .G(\pipeline/cu_pipeline/N113 ), 
        .D(\pipeline/cu_pipeline/N89 ), .Q(\pipeline/EXE_controls_in_IDEX[7] )
         );
  DLH_X1 \pipeline/cu_pipeline/Mem_to_reg_reg  ( .G(
        \pipeline/cu_pipeline/N107 ), .D(\pipeline/cu_pipeline/N108 ), .Q(
        \pipeline/WB_controls_in_IDEX[0] ) );
  DLL_X1 \pipeline/cu_pipeline/ALU_OPCODE_reg[1]  ( .D(
        \pipeline/cu_pipeline/N102 ), .GN(n13281), .Q(
        \pipeline/EXE_controls_in_IDEX[2] ) );
  DLH_X1 \pipeline/cu_pipeline/Alu_src_reg  ( .G(\pipeline/cu_pipeline/N112 ), 
        .D(\pipeline/cu_pipeline/N88 ), .Q(\pipeline/EXE_controls_in_IDEX[0] )
         );
  DLH_X1 \pipeline/cu_pipeline/isSigned_reg  ( .G(\pipeline/cu_pipeline/N109 ), 
        .D(\pipeline/cu_pipeline/N110 ), .Q(\pipeline/EXE_controls_in_IDEX[8] ) );
  DLL_X1 \pipeline/cu_pipeline/ALU_OPCODE_reg[4]  ( .D(
        \pipeline/cu_pipeline/N105 ), .GN(n13281), .Q(
        \pipeline/EXE_controls_in_IDEX[5] ) );
  DLH_X1 \pipeline/cu_hazard/stall_reg  ( .G(\pipeline/cu_hazard/N39 ), .D(
        \pipeline/cu_hazard/N40 ), .Q(\pipeline/stall ) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_tri_enable_reg[31]  ( .D(n3956), .CK(
        Clk), .RN(n17705), .Q(\pipeline/stageF/PC_reg/N0 ), .QN(n17379) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_tri_enable_reg[29]  ( .D(n3955), .CK(
        Clk), .RN(n17704), .Q(\pipeline/stageF/PC_reg/N2 ), .QN(n17494) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_tri_enable_reg[27]  ( .D(n3954), .CK(
        Clk), .RN(n17702), .Q(\pipeline/stageF/PC_reg/N4 ), .QN(n17493) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_tri_enable_reg[25]  ( .D(n3953), .CK(
        Clk), .RN(n17705), .Q(\pipeline/stageF/PC_reg/N6 ), .QN(n17492) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_tri_enable_reg[23]  ( .D(n3952), .CK(
        Clk), .RN(n17705), .Q(\pipeline/stageF/PC_reg/N8 ), .QN(n17491) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_tri_enable_reg[21]  ( .D(n3951), .CK(
        Clk), .RN(n17703), .Q(\pipeline/stageF/PC_reg/N10 ), .QN(n17490) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_tri_enable_reg[19]  ( .D(n3950), .CK(
        Clk), .RN(n17701), .Q(\pipeline/stageF/PC_reg/N12 ), .QN(n17489) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_tri_enable_reg[17]  ( .D(n3949), .CK(
        Clk), .RN(n17705), .Q(\pipeline/stageF/PC_reg/N14 ), .QN(n17488) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_tri_enable_reg[15]  ( .D(n3948), .CK(
        Clk), .RN(n17704), .Q(\pipeline/stageF/PC_reg/N16 ), .QN(n17487) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_tri_enable_reg[13]  ( .D(n3947), .CK(
        Clk), .RN(n17704), .Q(\pipeline/stageF/PC_reg/N18 ), .QN(n17486) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_tri_enable_reg[11]  ( .D(n3946), .CK(
        Clk), .RN(n17705), .Q(\pipeline/stageF/PC_reg/N20 ), .QN(n17485) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_tri_enable_reg[9]  ( .D(n3945), .CK(
        Clk), .RN(n17705), .Q(\pipeline/stageF/PC_reg/N22 ), .QN(n17378) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_tri_enable_reg[7]  ( .D(n3944), .CK(
        Clk), .RN(n17704), .Q(\pipeline/stageF/PC_reg/N24 ), .QN(n17484) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_tri_enable_reg[5]  ( .D(n3943), .CK(
        Clk), .RN(n17705), .Q(\pipeline/stageF/PC_reg/N26 ), .QN(n17483) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_tri_enable_reg[3]  ( .D(n3942), .CK(
        Clk), .RN(n17704), .Q(\pipeline/stageF/PC_reg/N28 ), .QN(n17482) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_tri_enable_reg[1]  ( .D(n3941), .CK(
        Clk), .RN(n17705), .Q(\pipeline/stageF/PC_reg/N30 ), .QN(n17377) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_tri_enable_reg[0]  ( .D(n3940), .CK(
        Clk), .RN(n17705), .Q(\pipeline/stageF/PC_reg/N31 ), .QN(n17376) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_tri_enable_reg[2]  ( .D(n3939), .CK(
        Clk), .RN(n17704), .Q(\pipeline/stageF/PC_reg/N29 ), .QN(n17481) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_tri_enable_reg[4]  ( .D(n3938), .CK(
        Clk), .RN(n17705), .Q(\pipeline/stageF/PC_reg/N27 ), .QN(n17480) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_tri_enable_reg[6]  ( .D(n3937), .CK(
        Clk), .RN(n17704), .Q(\pipeline/stageF/PC_reg/N25 ), .QN(n17479) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_tri_enable_reg[8]  ( .D(n3936), .CK(
        Clk), .RN(n17705), .Q(\pipeline/stageF/PC_reg/N23 ), .QN(n17478) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_tri_enable_reg[10]  ( .D(n3935), .CK(
        Clk), .RN(n17705), .Q(\pipeline/stageF/PC_reg/N21 ), .QN(n17375) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_tri_enable_reg[12]  ( .D(n3934), .CK(
        Clk), .RN(n17703), .Q(\pipeline/stageF/PC_reg/N19 ), .QN(n17477) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_tri_enable_reg[14]  ( .D(n3933), .CK(
        Clk), .RN(n17702), .Q(\pipeline/stageF/PC_reg/N17 ), .QN(n17476) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_tri_enable_reg[16]  ( .D(n3932), .CK(
        Clk), .RN(n17705), .Q(\pipeline/stageF/PC_reg/N15 ), .QN(n17475) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_tri_enable_reg[18]  ( .D(n3931), .CK(
        Clk), .RN(n17704), .Q(\pipeline/stageF/PC_reg/N13 ), .QN(n17474) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_tri_enable_reg[20]  ( .D(n3930), .CK(
        Clk), .RN(n17701), .Q(\pipeline/stageF/PC_reg/N11 ), .QN(n17473) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_tri_enable_reg[22]  ( .D(n3929), .CK(
        Clk), .RN(n17705), .Q(\pipeline/stageF/PC_reg/N9 ), .QN(n17374) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_tri_enable_reg[24]  ( .D(n3928), .CK(
        Clk), .RN(n17704), .Q(\pipeline/stageF/PC_reg/N7 ), .QN(n17472) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_tri_enable_reg[26]  ( .D(n3927), .CK(
        Clk), .RN(n17705), .Q(\pipeline/stageF/PC_reg/N5 ), .QN(n17373) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_tri_enable_reg[28]  ( .D(n3926), .CK(
        Clk), .RN(n17705), .Q(\pipeline/stageF/PC_reg/N3 ), .QN(n17372) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_tri_enable_reg[30]  ( .D(n3925), .CK(
        Clk), .RN(n17705), .Q(\pipeline/stageF/PC_reg/N1 ), .QN(n17371) );
  DFF_X1 \pipeline/IDEX_Stage/MEM_controls_out_IDEX_reg[1]  ( .D(
        \pipeline/IDEX_Stage/N92 ), .CK(Clk), .Q(
        \pipeline/MEM_controls_in_EXMEM[1] ) );
  DFF_X1 \pipeline/EXMEM_stage/MEM_controls_out_EXMEM_reg[1]  ( .D(
        \pipeline/EXMEM_stage/N6 ), .CK(Clk), .Q(
        \pipeline/MEM_controls_in_MEM[1] ), .QN(n17019) );
  DFF_X1 \pipeline/IDEX_Stage/MEM_controls_out_IDEX_reg[0]  ( .D(
        \pipeline/IDEX_Stage/N91 ), .CK(Clk), .Q(n13942), .QN(n17447) );
  DFF_X1 \pipeline/EXMEM_stage/MEM_controls_out_EXMEM_reg[0]  ( .D(
        \pipeline/EXMEM_stage/N5 ), .CK(Clk), .QN(n17020) );
  DLL_X1 \pipeline/stageM/read_notWrite_reg  ( .D(
        \pipeline/MEM_controls_in_MEM[1] ), .GN(n17155), .Q(read_notWrite) );
  DLL_X1 \DataMem/Dataout_tri_enable_reg[31]  ( .D(n17155), .GN(n17098), .Q(
        \DataMem/N0 ) );
  DLL_X1 \DataMem/Dataout_tri_enable_reg[29]  ( .D(n12766), .GN(n17098), .Q(
        \DataMem/N2 ) );
  DLL_X1 \DataMem/Dataout_tri_enable_reg[27]  ( .D(n12766), .GN(n17098), .Q(
        \DataMem/N4 ) );
  DLL_X1 \DataMem/Dataout_tri_enable_reg[25]  ( .D(n17155), .GN(n17098), .Q(
        \DataMem/N6 ) );
  DLL_X1 \DataMem/Dataout_tri_enable_reg[23]  ( .D(n17155), .GN(n13055), .Q(
        \DataMem/N8 ) );
  DLL_X1 \DataMem/Dataout_tri_enable_reg[21]  ( .D(n12766), .GN(n17098), .Q(
        \DataMem/N10 ) );
  DLL_X1 \DataMem/Dataout_tri_enable_reg[19]  ( .D(n17155), .GN(n17098), .Q(
        \DataMem/N12 ) );
  DLL_X1 \DataMem/Dataout_tri_enable_reg[17]  ( .D(n12766), .GN(n17098), .Q(
        \DataMem/N14 ) );
  DLL_X1 \DataMem/Dataout_tri_enable_reg[15]  ( .D(n12766), .GN(n17098), .Q(
        \DataMem/N16 ) );
  DLL_X1 \DataMem/Dataout_tri_enable_reg[13]  ( .D(n17155), .GN(n17098), .Q(
        \DataMem/N18 ) );
  DLL_X1 \DataMem/Dataout_tri_enable_reg[11]  ( .D(n12766), .GN(n17098), .Q(
        \DataMem/N20 ) );
  DLL_X1 \DataMem/Dataout_tri_enable_reg[9]  ( .D(n17155), .GN(n17098), .Q(
        \DataMem/N22 ) );
  DLL_X1 \DataMem/Dataout_tri_enable_reg[7]  ( .D(n17155), .GN(n17098), .Q(
        \DataMem/N24 ) );
  DLL_X1 \DataMem/Dataout_tri_enable_reg[5]  ( .D(n12766), .GN(n17098), .Q(
        \DataMem/N26 ) );
  DLL_X1 \DataMem/Dataout_tri_enable_reg[3]  ( .D(n17155), .GN(n17098), .Q(
        \DataMem/N28 ) );
  DLL_X1 \DataMem/Dataout_tri_enable_reg[1]  ( .D(n12766), .GN(n17098), .Q(
        \DataMem/N30 ) );
  DLL_X1 \DataMem/Dataout_tri_enable_reg[0]  ( .D(n17155), .GN(n17098), .Q(
        \DataMem/N31 ) );
  DLL_X1 \DataMem/Dataout_tri_enable_reg[2]  ( .D(n12766), .GN(n17098), .Q(
        \DataMem/N29 ) );
  DLL_X1 \DataMem/Dataout_tri_enable_reg[4]  ( .D(n17155), .GN(n17098), .Q(
        \DataMem/N27 ) );
  DLL_X1 \DataMem/Dataout_tri_enable_reg[6]  ( .D(n17155), .GN(n17098), .Q(
        \DataMem/N25 ) );
  DLL_X1 \DataMem/Dataout_tri_enable_reg[8]  ( .D(n12766), .GN(n17098), .Q(
        \DataMem/N23 ) );
  DLL_X1 \DataMem/Dataout_tri_enable_reg[10]  ( .D(n17155), .GN(n17098), .Q(
        \DataMem/N21 ) );
  DLL_X1 \DataMem/Dataout_tri_enable_reg[12]  ( .D(n12766), .GN(n17098), .Q(
        \DataMem/N19 ) );
  DLL_X1 \DataMem/Dataout_tri_enable_reg[14]  ( .D(n12766), .GN(n17098), .Q(
        \DataMem/N17 ) );
  DLL_X1 \DataMem/Dataout_tri_enable_reg[16]  ( .D(n17155), .GN(n17098), .Q(
        \DataMem/N15 ) );
  DLL_X1 \DataMem/Dataout_tri_enable_reg[18]  ( .D(n17155), .GN(n17098), .Q(
        \DataMem/N13 ) );
  DLL_X1 \DataMem/Dataout_tri_enable_reg[20]  ( .D(n17155), .GN(n17098), .Q(
        \DataMem/N11 ) );
  DLL_X1 \DataMem/Dataout_tri_enable_reg[22]  ( .D(n17155), .GN(n17098), .Q(
        \DataMem/N9 ) );
  DLL_X1 \DataMem/Dataout_tri_enable_reg[24]  ( .D(n12766), .GN(n17098), .Q(
        \DataMem/N7 ) );
  DLL_X1 \DataMem/Dataout_tri_enable_reg[26]  ( .D(n12766), .GN(n17098), .Q(
        \DataMem/N5 ) );
  DLL_X1 \DataMem/Dataout_tri_enable_reg[28]  ( .D(n12766), .GN(n17098), .Q(
        \DataMem/N3 ) );
  DLL_X1 \DataMem/Dataout_tri_enable_reg[30]  ( .D(n17155), .GN(n17098), .Q(
        \DataMem/N1 ) );
  DFF_X1 \pipeline/IDEX_Stage/WB_controls_out_IDEX_reg[1]  ( .D(
        \pipeline/IDEX_Stage/N90 ), .CK(Clk), .Q(
        \pipeline/WB_controls_in_EXMEM[1] ), .QN(n17449) );
  DFF_X1 \pipeline/EXMEM_stage/WB_controls_out_EXMEM_reg[1]  ( .D(
        \pipeline/EXMEM_stage/N4 ), .CK(Clk), .Q(
        \pipeline/WB_controls_in_MEMWB[1] ), .QN(n17387) );
  DFF_X1 \pipeline/MEMWB_Stage/writeback_reg  ( .D(\pipeline/MEMWB_Stage/N10 ), 
        .CK(Clk), .QN(n13940) );
  DFF_X1 \pipeline/IDEX_Stage/EXE_controls_out_IDEX_reg[8]  ( .D(
        \pipeline/IDEX_Stage/N101 ), .CK(Clk), .Q(n13939) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_reg[31]  ( .D(n3924), .CK(Clk), .RN(
        n17705), .Q(n13938), .QN(n7676) );
  DFF_X1 \pipeline/IFID_stage/PC_out_IFID_reg[31]  ( .D(n3923), .CK(Clk), .Q(
        n13937), .QN(n17527) );
  DFF_X1 \pipeline/IDEX_Stage/EXE_controls_out_IDEX_reg[6]  ( .D(
        \pipeline/IDEX_Stage/N99 ), .CK(Clk), .Q(
        \pipeline/EXE_controls_in_EXEcute [6]), .QN(n17421) );
  DFF_X1 \pipeline/IDEX_Stage/EXE_controls_out_IDEX_reg[5]  ( .D(
        \pipeline/IDEX_Stage/N98 ), .CK(Clk), .Q(
        \pipeline/EXE_controls_in_EXEcute [5]) );
  DFF_X1 \pipeline/IDEX_Stage/EXE_controls_out_IDEX_reg[4]  ( .D(
        \pipeline/IDEX_Stage/N97 ), .CK(Clk), .Q(
        \pipeline/EXE_controls_in_EXEcute [4]) );
  DFF_X1 \pipeline/IDEX_Stage/EXE_controls_out_IDEX_reg[3]  ( .D(
        \pipeline/IDEX_Stage/N96 ), .CK(Clk), .Q(
        \pipeline/EXE_controls_in_EXEcute [3]), .QN(n17411) );
  DFF_X1 \pipeline/IDEX_Stage/EXE_controls_out_IDEX_reg[2]  ( .D(
        \pipeline/IDEX_Stage/N95 ), .CK(Clk), .Q(
        \pipeline/EXE_controls_in_EXEcute [2]), .QN(n17405) );
  DFF_X1 \pipeline/IDEX_Stage/WB_controls_out_IDEX_reg[0]  ( .D(
        \pipeline/IDEX_Stage/N89 ), .CK(Clk), .Q(n13936) );
  DFF_X1 \pipeline/EXMEM_stage/WB_controls_out_EXMEM_reg[0]  ( .D(
        \pipeline/EXMEM_stage/N3 ), .CK(Clk), .Q(
        \pipeline/WB_controls_in_MEMWB[0] ) );
  DFF_X1 \pipeline/IDEX_Stage/RegDst_2_Addr_out_IDEX_reg[4]  ( .D(
        \pipeline/IDEX_Stage/N217 ), .CK(Clk), .Q(n13934) );
  DFF_X1 \pipeline/IDEX_Stage/RegDst_2_Addr_out_IDEX_reg[3]  ( .D(
        \pipeline/IDEX_Stage/N216 ), .CK(Clk), .Q(n13933) );
  DFF_X1 \pipeline/IDEX_Stage/RegDst_2_Addr_out_IDEX_reg[2]  ( .D(
        \pipeline/IDEX_Stage/N215 ), .CK(Clk), .Q(n13932) );
  DFF_X1 \pipeline/IDEX_Stage/RegDst_2_Addr_out_IDEX_reg[1]  ( .D(
        \pipeline/IDEX_Stage/N214 ), .CK(Clk), .Q(n13931) );
  DFF_X1 \pipeline/IDEX_Stage/RegDst_2_Addr_out_IDEX_reg[0]  ( .D(
        \pipeline/IDEX_Stage/N213 ), .CK(Clk), .Q(n13930) );
  DFF_X1 \pipeline/IDEX_Stage/RegDst_1_Addr_out_IDEX_reg[4]  ( .D(
        \pipeline/IDEX_Stage/N212 ), .CK(Clk), .Q(n13929) );
  DFF_X1 \pipeline/IDEX_Stage/RegDst_1_Addr_out_IDEX_reg[3]  ( .D(
        \pipeline/IDEX_Stage/N211 ), .CK(Clk), .Q(n13928) );
  DFF_X1 \pipeline/IDEX_Stage/RegDst_1_Addr_out_IDEX_reg[2]  ( .D(
        \pipeline/IDEX_Stage/N210 ), .CK(Clk), .Q(n13927) );
  DFF_X1 \pipeline/IDEX_Stage/RegDst_1_Addr_out_IDEX_reg[1]  ( .D(
        \pipeline/IDEX_Stage/N209 ), .CK(Clk), .Q(n13926) );
  DFF_X1 \pipeline/IDEX_Stage/RegDst_1_Addr_out_IDEX_reg[0]  ( .D(
        \pipeline/IDEX_Stage/N208 ), .CK(Clk), .Q(n13925) );
  DFF_X1 \pipeline/IDEX_Stage/Immediate_out_IDEX_reg[2]  ( .D(
        \pipeline/IDEX_Stage/N168 ), .CK(Clk), .Q(
        \pipeline/immediate_to_exe [2]) );
  DFF_X1 \pipeline/IDEX_Stage/Reg2_Addr_out_IDEX_reg[3]  ( .D(
        \pipeline/IDEX_Stage/N206 ), .CK(Clk), .Q(
        \pipeline/Reg2_Addr_to_exe [3]) );
  DFF_X1 \pipeline/IDEX_Stage/Reg2_Addr_out_IDEX_reg[2]  ( .D(
        \pipeline/IDEX_Stage/N205 ), .CK(Clk), .Q(
        \pipeline/Reg2_Addr_to_exe [2]), .QN(n17403) );
  DFF_X1 \pipeline/IDEX_Stage/Reg2_Addr_out_IDEX_reg[0]  ( .D(
        \pipeline/IDEX_Stage/N203 ), .CK(Clk), .Q(
        \pipeline/Reg2_Addr_to_exe [0]) );
  DFF_X1 \pipeline/IDEX_Stage/Reg1_Addr_out_IDEX_reg[4]  ( .D(
        \pipeline/IDEX_Stage/N202 ), .CK(Clk), .Q(
        \pipeline/Reg1_Addr_to_exe [4]), .QN(n17399) );
  DFF_X1 \pipeline/IDEX_Stage/Reg1_Addr_out_IDEX_reg[3]  ( .D(
        \pipeline/IDEX_Stage/N201 ), .CK(Clk), .Q(
        \pipeline/Reg1_Addr_to_exe [3]) );
  DFF_X1 \pipeline/IDEX_Stage/Reg1_Addr_out_IDEX_reg[2]  ( .D(
        \pipeline/IDEX_Stage/N200 ), .CK(Clk), .Q(
        \pipeline/Reg1_Addr_to_exe [2]), .QN(n17401) );
  DFF_X1 \pipeline/IDEX_Stage/Reg1_Addr_out_IDEX_reg[1]  ( .D(
        \pipeline/IDEX_Stage/N199 ), .CK(Clk), .Q(
        \pipeline/Reg1_Addr_to_exe [1]) );
  DFF_X1 \pipeline/IDEX_Stage/Immediate_out_IDEX_reg[15]  ( .D(
        \pipeline/IDEX_Stage/N181 ), .CK(Clk), .Q(
        \pipeline/immediate_to_exe [15]) );
  DFF_X1 \pipeline/IDEX_Stage/Immediate_out_IDEX_reg[13]  ( .D(
        \pipeline/IDEX_Stage/N179 ), .CK(Clk), .Q(
        \pipeline/immediate_to_exe [13]) );
  DFF_X1 \pipeline/IDEX_Stage/Immediate_out_IDEX_reg[12]  ( .D(
        \pipeline/IDEX_Stage/N178 ), .CK(Clk), .Q(
        \pipeline/immediate_to_exe [12]) );
  DFF_X1 \pipeline/IDEX_Stage/Immediate_out_IDEX_reg[11]  ( .D(
        \pipeline/IDEX_Stage/N177 ), .CK(Clk), .Q(
        \pipeline/immediate_to_exe [11]) );
  DFF_X1 \pipeline/IDEX_Stage/Immediate_out_IDEX_reg[9]  ( .D(
        \pipeline/IDEX_Stage/N175 ), .CK(Clk), .Q(
        \pipeline/immediate_to_exe [9]) );
  DFF_X1 \pipeline/IDEX_Stage/Immediate_out_IDEX_reg[8]  ( .D(
        \pipeline/IDEX_Stage/N174 ), .CK(Clk), .Q(
        \pipeline/immediate_to_exe [8]) );
  DFF_X1 \pipeline/IDEX_Stage/Immediate_out_IDEX_reg[7]  ( .D(
        \pipeline/IDEX_Stage/N173 ), .CK(Clk), .Q(
        \pipeline/immediate_to_exe [7]) );
  DFF_X1 \pipeline/IDEX_Stage/Immediate_out_IDEX_reg[31]  ( .D(
        \pipeline/IDEX_Stage/N197 ), .CK(Clk), .Q(
        \pipeline/immediate_to_exe [31]) );
  DFF_X1 \pipeline/IDEX_Stage/Immediate_out_IDEX_reg[29]  ( .D(
        \pipeline/IDEX_Stage/N197 ), .CK(Clk), .Q(
        \pipeline/immediate_to_exe [29]) );
  DFF_X1 \pipeline/IDEX_Stage/Immediate_out_IDEX_reg[27]  ( .D(
        \pipeline/IDEX_Stage/N197 ), .CK(Clk), .Q(
        \pipeline/immediate_to_exe [27]) );
  DFF_X1 \pipeline/IDEX_Stage/Immediate_out_IDEX_reg[25]  ( .D(
        \pipeline/IDEX_Stage/N197 ), .CK(Clk), .Q(
        \pipeline/immediate_to_exe [25]) );
  DFF_X1 \pipeline/IDEX_Stage/Immediate_out_IDEX_reg[23]  ( .D(
        \pipeline/IDEX_Stage/N197 ), .CK(Clk), .Q(
        \pipeline/immediate_to_exe [23]) );
  DFF_X1 \pipeline/IDEX_Stage/Immediate_out_IDEX_reg[21]  ( .D(
        \pipeline/IDEX_Stage/N197 ), .CK(Clk), .Q(
        \pipeline/immediate_to_exe [21]) );
  DFF_X1 \pipeline/IDEX_Stage/Immediate_out_IDEX_reg[19]  ( .D(
        \pipeline/IDEX_Stage/N197 ), .CK(Clk), .Q(
        \pipeline/immediate_to_exe [19]) );
  DFF_X1 \pipeline/IDEX_Stage/Immediate_out_IDEX_reg[17]  ( .D(
        \pipeline/IDEX_Stage/N197 ), .CK(Clk), .Q(
        \pipeline/immediate_to_exe [17]) );
  DFF_X1 \pipeline/IDEX_Stage/Immediate_out_IDEX_reg[16]  ( .D(
        \pipeline/IDEX_Stage/N197 ), .CK(Clk), .Q(
        \pipeline/immediate_to_exe [16]) );
  DFF_X1 \pipeline/IDEX_Stage/Immediate_out_IDEX_reg[18]  ( .D(
        \pipeline/IDEX_Stage/N197 ), .CK(Clk), .Q(
        \pipeline/immediate_to_exe [18]) );
  DFF_X1 \pipeline/IDEX_Stage/Immediate_out_IDEX_reg[20]  ( .D(
        \pipeline/IDEX_Stage/N197 ), .CK(Clk), .Q(
        \pipeline/immediate_to_exe [20]) );
  DFF_X1 \pipeline/IDEX_Stage/Immediate_out_IDEX_reg[22]  ( .D(
        \pipeline/IDEX_Stage/N197 ), .CK(Clk), .Q(
        \pipeline/immediate_to_exe [22]) );
  DFF_X1 \pipeline/IDEX_Stage/Immediate_out_IDEX_reg[24]  ( .D(
        \pipeline/IDEX_Stage/N197 ), .CK(Clk), .Q(
        \pipeline/immediate_to_exe [24]) );
  DFF_X1 \pipeline/IDEX_Stage/Immediate_out_IDEX_reg[26]  ( .D(
        \pipeline/IDEX_Stage/N197 ), .CK(Clk), .Q(
        \pipeline/immediate_to_exe [26]) );
  DFF_X1 \pipeline/IDEX_Stage/Immediate_out_IDEX_reg[28]  ( .D(
        \pipeline/IDEX_Stage/N197 ), .CK(Clk), .Q(
        \pipeline/immediate_to_exe [28]) );
  DFF_X1 \pipeline/IDEX_Stage/Immediate_out_IDEX_reg[30]  ( .D(
        \pipeline/IDEX_Stage/N197 ), .CK(Clk), .Q(
        \pipeline/immediate_to_exe [30]) );
  DFF_X1 \pipeline/IDEX_Stage/Immediate_out_IDEX_reg[10]  ( .D(
        \pipeline/IDEX_Stage/N176 ), .CK(Clk), .Q(
        \pipeline/immediate_to_exe [10]) );
  DFF_X1 \pipeline/IDEX_Stage/Immediate_out_IDEX_reg[6]  ( .D(
        \pipeline/IDEX_Stage/N172 ), .CK(Clk), .Q(
        \pipeline/immediate_to_exe [6]) );
  DFF_X1 \pipeline/IDEX_Stage/Immediate_out_IDEX_reg[5]  ( .D(
        \pipeline/IDEX_Stage/N171 ), .CK(Clk), .Q(
        \pipeline/immediate_to_exe [5]) );
  DFF_X1 \pipeline/IDEX_Stage/Immediate_out_IDEX_reg[4]  ( .D(
        \pipeline/IDEX_Stage/N170 ), .CK(Clk), .Q(
        \pipeline/immediate_to_exe [4]) );
  DFF_X1 \pipeline/IDEX_Stage/Immediate_out_IDEX_reg[3]  ( .D(
        \pipeline/IDEX_Stage/N169 ), .CK(Clk), .Q(
        \pipeline/immediate_to_exe [3]) );
  DFF_X1 \pipeline/IDEX_Stage/Immediate_out_IDEX_reg[1]  ( .D(
        \pipeline/IDEX_Stage/N167 ), .CK(Clk), .Q(
        \pipeline/immediate_to_exe [1]) );
  DFF_X1 \pipeline/IDEX_Stage/Immediate_out_IDEX_reg[0]  ( .D(
        \pipeline/IDEX_Stage/N166 ), .CK(Clk), .QN(n17400) );
  DFF_X1 \pipeline/IDEX_Stage/EXE_controls_out_IDEX_reg[7]  ( .D(
        \pipeline/IDEX_Stage/N100 ), .CK(Clk), .Q(
        \pipeline/EXE_controls_in_EXEcute [7]), .QN(n17430) );
  DFF_X1 \pipeline/MEMWB_Stage/RegDst_Addr_out_MEMWB_reg[3]  ( .D(
        \pipeline/MEMWB_Stage/N46 ), .CK(Clk), .Q(\pipeline/RegDst_to_WB[3] ), 
        .QN(n17385) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[2][31]  ( .G(n13169), .D(n13268), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[2][31] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[2][29]  ( .G(n17707), .D(n13262), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[2][29] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[2][27]  ( .G(n13169), .D(n13256), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[2][27] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[2][25]  ( .G(n17707), .D(n13250), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[2][25] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[2][23]  ( .G(n17707), .D(n13244), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[2][23] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[2][21]  ( .G(n13169), .D(n13238), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[2][21] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[2][19]  ( .G(n17707), .D(n13232), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[2][19] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[2][17]  ( .G(n13169), .D(n13226), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[2][17] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[2][15]  ( .G(n17707), .D(n13220), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[2][15] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[2][13]  ( .G(n13169), .D(n13214), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[2][13] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[2][0]  ( .G(n17707), .D(n13175), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[2][0] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[2][8]  ( .G(n17707), .D(n13199), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[2][8] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[2][14]  ( .G(n13169), .D(n13217), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[2][14] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[2][16]  ( .G(n17707), .D(n13223), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[2][16] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[2][18]  ( .G(n17707), .D(n13229), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[2][18] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[2][20]  ( .G(n13169), .D(n13235), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[2][20] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[2][22]  ( .G(n13169), .D(n13241), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[2][22] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[2][24]  ( .G(n13169), .D(n13247), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[2][24] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[2][26]  ( .G(n13169), .D(n13253), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[2][26] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[2][28]  ( .G(n13169), .D(n13259), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[2][28] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[2][30]  ( .G(n17707), .D(n13265), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[2][30] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[3][31]  ( .G(n17708), .D(n13268), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[3][31] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[3][29]  ( .G(n17708), .D(n13262), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[3][29] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[3][27]  ( .G(n13166), .D(n13256), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[3][27] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[3][25]  ( .G(n17708), .D(n13250), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[3][25] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[3][23]  ( .G(n13166), .D(n13244), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[3][23] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[3][21]  ( .G(n13166), .D(n13238), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[3][21] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[3][19]  ( .G(n17708), .D(n13232), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[3][19] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[3][17]  ( .G(n13166), .D(n13226), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[3][17] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[3][15]  ( .G(n17708), .D(n13220), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[3][15] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[3][13]  ( .G(n13166), .D(n13214), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[3][13] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[3][0]  ( .G(n17708), .D(n13175), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[3][0] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[3][8]  ( .G(n17708), .D(n13199), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[3][8] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[3][14]  ( .G(n13166), .D(n13217), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[3][14] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[3][16]  ( .G(n17708), .D(n13223), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[3][16] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[3][18]  ( .G(n17708), .D(n13229), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[3][18] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[3][20]  ( .G(n13166), .D(n13235), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[3][20] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[3][22]  ( .G(n13166), .D(n13241), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[3][22] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[3][24]  ( .G(n13166), .D(n13247), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[3][24] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[3][26]  ( .G(n13166), .D(n13253), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[3][26] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[3][28]  ( .G(n13166), .D(n13259), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[3][28] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[3][30]  ( .G(n17708), .D(n13265), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[3][30] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[4][31]  ( .G(n13163), .D(n13268), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[4][31] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[4][29]  ( .G(n17709), .D(n13262), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[4][29] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[4][27]  ( .G(n13163), .D(n13256), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[4][27] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[4][25]  ( .G(n17709), .D(n13250), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[4][25] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[4][23]  ( .G(n17709), .D(n13244), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[4][23] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[4][21]  ( .G(n13163), .D(n13238), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[4][21] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[4][19]  ( .G(n17709), .D(n13232), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[4][19] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[4][17]  ( .G(n13163), .D(n13226), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[4][17] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[4][15]  ( .G(n17709), .D(n13220), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[4][15] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[4][13]  ( .G(n13163), .D(n13214), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[4][13] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[4][0]  ( .G(n17709), .D(n13175), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[4][0] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[4][8]  ( .G(n17709), .D(n13199), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[4][8] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[4][14]  ( .G(n13163), .D(n13217), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[4][14] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[4][16]  ( .G(n17709), .D(n13223), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[4][16] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[4][18]  ( .G(n17709), .D(n13229), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[4][18] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[4][20]  ( .G(n13163), .D(n13235), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[4][20] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[4][22]  ( .G(n13163), .D(n13241), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[4][22] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[4][24]  ( .G(n13163), .D(n13247), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[4][24] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[4][26]  ( .G(n13163), .D(n13253), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[4][26] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[4][28]  ( .G(n13163), .D(n13259), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[4][28] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[4][30]  ( .G(n17709), .D(n13265), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[4][30] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[5][31]  ( .G(n13160), .D(n13268), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[5][31] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[5][29]  ( .G(n17710), .D(n13262), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[5][29] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[5][27]  ( .G(n13160), .D(n13256), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[5][27] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[5][25]  ( .G(n17710), .D(n13250), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[5][25] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[5][23]  ( .G(n17710), .D(n13244), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[5][23] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[5][21]  ( .G(n13160), .D(n13238), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[5][21] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[5][19]  ( .G(n17710), .D(n13232), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[5][19] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[5][17]  ( .G(n13160), .D(n13226), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[5][17] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[5][15]  ( .G(n17710), .D(n13220), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[5][15] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[5][13]  ( .G(n13160), .D(n13214), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[5][13] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[5][0]  ( .G(n17710), .D(n13175), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[5][0] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[5][8]  ( .G(n17710), .D(n13199), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[5][8] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[5][14]  ( .G(n13160), .D(n13217), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[5][14] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[5][16]  ( .G(n17710), .D(n13223), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[5][16] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[5][18]  ( .G(n17710), .D(n13229), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[5][18] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[5][20]  ( .G(n13160), .D(n13235), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[5][20] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[5][22]  ( .G(n13160), .D(n13241), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[5][22] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[5][24]  ( .G(n13160), .D(n13247), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[5][24] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[5][26]  ( .G(n13160), .D(n13253), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[5][26] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[5][28]  ( .G(n13160), .D(n13259), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[5][28] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[5][30]  ( .G(n17710), .D(n13265), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[5][30] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[6][31]  ( .G(n13157), .D(n13268), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[6][31] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[6][29]  ( .G(n17711), .D(n13262), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[6][29] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[6][27]  ( .G(n13157), .D(n13256), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[6][27] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[6][25]  ( .G(n17711), .D(n13250), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[6][25] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[6][23]  ( .G(n17711), .D(n13244), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[6][23] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[6][21]  ( .G(n13157), .D(n13238), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[6][21] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[6][19]  ( .G(n17711), .D(n13232), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[6][19] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[6][17]  ( .G(n13157), .D(n13226), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[6][17] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[6][15]  ( .G(n17711), .D(n13220), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[6][15] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[6][13]  ( .G(n13157), .D(n13214), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[6][13] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[6][0]  ( .G(n17711), .D(n13175), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[6][0] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[6][8]  ( .G(n17711), .D(n13199), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[6][8] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[6][14]  ( .G(n13157), .D(n13217), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[6][14] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[6][16]  ( .G(n17711), .D(n13223), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[6][16] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[6][18]  ( .G(n17711), .D(n13229), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[6][18] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[6][20]  ( .G(n13157), .D(n13235), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[6][20] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[6][22]  ( .G(n13157), .D(n13241), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[6][22] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[6][24]  ( .G(n13157), .D(n13247), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[6][24] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[6][26]  ( .G(n13157), .D(n13253), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[6][26] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[6][28]  ( .G(n13157), .D(n13259), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[6][28] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[6][30]  ( .G(n17711), .D(n13265), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[6][30] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[7][31]  ( .G(n13154), .D(n13268), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[7][31] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[7][29]  ( .G(n17712), .D(n13262), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[7][29] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[7][27]  ( .G(n13154), .D(n13256), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[7][27] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[7][25]  ( .G(n17712), .D(n13250), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[7][25] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[7][23]  ( .G(n17712), .D(n13244), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[7][23] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[7][21]  ( .G(n13154), .D(n13238), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[7][21] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[7][19]  ( .G(n17712), .D(n13232), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[7][19] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[7][17]  ( .G(n13154), .D(n13226), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[7][17] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[7][15]  ( .G(n17712), .D(n13220), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[7][15] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[7][13]  ( .G(n13154), .D(n13214), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[7][13] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[7][0]  ( .G(n17712), .D(n13175), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[7][0] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[7][8]  ( .G(n17712), .D(n13199), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[7][8] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[7][14]  ( .G(n13154), .D(n13217), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[7][14] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[7][16]  ( .G(n17712), .D(n13223), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[7][16] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[7][18]  ( .G(n17712), .D(n13229), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[7][18] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[7][20]  ( .G(n13154), .D(n13235), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[7][20] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[7][22]  ( .G(n13154), .D(n13241), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[7][22] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[7][24]  ( .G(n13154), .D(n13247), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[7][24] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[7][26]  ( .G(n13154), .D(n13253), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[7][26] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[7][28]  ( .G(n13154), .D(n13259), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[7][28] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[7][30]  ( .G(n17712), .D(n13265), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[7][30] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[8][31]  ( .G(n13151), .D(n13268), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[8][31] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[8][29]  ( .G(n17713), .D(n13262), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[8][29] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[8][27]  ( .G(n13151), .D(n13256), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[8][27] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[8][25]  ( .G(n17713), .D(n13250), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[8][25] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[8][23]  ( .G(n17713), .D(n13244), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[8][23] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[8][21]  ( .G(n13151), .D(n13238), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[8][21] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[8][19]  ( .G(n17713), .D(n13232), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[8][19] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[8][17]  ( .G(n13151), .D(n13226), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[8][17] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[8][15]  ( .G(n17713), .D(n13220), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[8][15] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[8][13]  ( .G(n13151), .D(n13214), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[8][13] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[8][0]  ( .G(n17713), .D(n13175), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[8][0] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[8][8]  ( .G(n17713), .D(n13199), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[8][8] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[8][14]  ( .G(n13151), .D(n13217), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[8][14] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[8][16]  ( .G(n17713), .D(n13223), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[8][16] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[8][18]  ( .G(n17713), .D(n13229), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[8][18] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[8][20]  ( .G(n13151), .D(n13235), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[8][20] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[8][22]  ( .G(n13151), .D(n13241), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[8][22] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[8][24]  ( .G(n13151), .D(n13247), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[8][24] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[8][26]  ( .G(n13151), .D(n13253), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[8][26] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[8][28]  ( .G(n13151), .D(n13259), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[8][28] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[8][30]  ( .G(n17713), .D(n13265), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[8][30] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[9][31]  ( .G(n13148), .D(n13268), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[9][31] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[9][29]  ( .G(n17714), .D(n13262), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[9][29] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[9][27]  ( .G(n13148), .D(n13256), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[9][27] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[9][25]  ( .G(n17714), .D(n13250), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[9][25] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[9][23]  ( .G(n17714), .D(n13244), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[9][23] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[9][21]  ( .G(n13148), .D(n13238), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[9][21] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[9][19]  ( .G(n17714), .D(n13232), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[9][19] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[9][17]  ( .G(n13148), .D(n13226), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[9][17] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[9][15]  ( .G(n17714), .D(n13220), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[9][15] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[9][13]  ( .G(n13148), .D(n13214), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[9][13] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[9][0]  ( .G(n17714), .D(n13175), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[9][0] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[9][8]  ( .G(n17714), .D(n13199), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[9][8] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[9][14]  ( .G(n13148), .D(n13217), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[9][14] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[9][16]  ( .G(n17714), .D(n13223), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[9][16] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[9][18]  ( .G(n17714), .D(n13229), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[9][18] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[9][20]  ( .G(n13148), .D(n13235), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[9][20] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[9][22]  ( .G(n13148), .D(n13241), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[9][22] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[9][24]  ( .G(n13148), .D(n13247), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[9][24] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[9][26]  ( .G(n13148), .D(n13253), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[9][26] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[9][28]  ( .G(n13148), .D(n13259), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[9][28] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[9][30]  ( .G(n17714), .D(n13265), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[9][30] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[10][31]  ( .G(n13145), .D(n13268), .Q(\pipeline/RegFile_DEC_WB/RegBank[10][31] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[10][29]  ( .G(n17715), .D(n13262), .Q(\pipeline/RegFile_DEC_WB/RegBank[10][29] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[10][27]  ( .G(n13145), .D(n13256), .Q(\pipeline/RegFile_DEC_WB/RegBank[10][27] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[10][25]  ( .G(n17715), .D(n13250), .Q(\pipeline/RegFile_DEC_WB/RegBank[10][25] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[10][23]  ( .G(n17715), .D(n13244), .Q(\pipeline/RegFile_DEC_WB/RegBank[10][23] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[10][21]  ( .G(n13145), .D(n13238), .Q(\pipeline/RegFile_DEC_WB/RegBank[10][21] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[10][19]  ( .G(n17715), .D(n13232), .Q(\pipeline/RegFile_DEC_WB/RegBank[10][19] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[10][17]  ( .G(n13145), .D(n13226), .Q(\pipeline/RegFile_DEC_WB/RegBank[10][17] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[10][15]  ( .G(n17715), .D(n13220), .Q(\pipeline/RegFile_DEC_WB/RegBank[10][15] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[10][13]  ( .G(n13145), .D(n13214), .Q(\pipeline/RegFile_DEC_WB/RegBank[10][13] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[10][0]  ( .G(n17715), .D(n13175), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[10][0] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[10][8]  ( .G(n17715), .D(n13199), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[10][8] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[10][14]  ( .G(n13145), .D(n13217), .Q(\pipeline/RegFile_DEC_WB/RegBank[10][14] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[10][16]  ( .G(n17715), .D(n13223), .Q(\pipeline/RegFile_DEC_WB/RegBank[10][16] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[10][18]  ( .G(n17715), .D(n13229), .Q(\pipeline/RegFile_DEC_WB/RegBank[10][18] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[10][20]  ( .G(n13145), .D(n13235), .Q(\pipeline/RegFile_DEC_WB/RegBank[10][20] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[10][22]  ( .G(n13145), .D(n13241), .Q(\pipeline/RegFile_DEC_WB/RegBank[10][22] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[10][24]  ( .G(n13145), .D(n13247), .Q(\pipeline/RegFile_DEC_WB/RegBank[10][24] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[10][26]  ( .G(n13145), .D(n13253), .Q(\pipeline/RegFile_DEC_WB/RegBank[10][26] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[10][28]  ( .G(n13145), .D(n13259), .Q(\pipeline/RegFile_DEC_WB/RegBank[10][28] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[10][30]  ( .G(n17715), .D(n13265), .Q(\pipeline/RegFile_DEC_WB/RegBank[10][30] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[11][31]  ( .G(n13142), .D(n13268), .Q(\pipeline/RegFile_DEC_WB/RegBank[11][31] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[11][29]  ( .G(n17716), .D(n13262), .Q(\pipeline/RegFile_DEC_WB/RegBank[11][29] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[11][27]  ( .G(n13142), .D(n13256), .Q(\pipeline/RegFile_DEC_WB/RegBank[11][27] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[11][25]  ( .G(n17716), .D(n13250), .Q(\pipeline/RegFile_DEC_WB/RegBank[11][25] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[11][23]  ( .G(n17716), .D(n13244), .Q(\pipeline/RegFile_DEC_WB/RegBank[11][23] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[11][21]  ( .G(n13142), .D(n13238), .Q(\pipeline/RegFile_DEC_WB/RegBank[11][21] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[11][19]  ( .G(n17716), .D(n13232), .Q(\pipeline/RegFile_DEC_WB/RegBank[11][19] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[11][17]  ( .G(n13142), .D(n13226), .Q(\pipeline/RegFile_DEC_WB/RegBank[11][17] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[11][15]  ( .G(n17716), .D(n13220), .Q(\pipeline/RegFile_DEC_WB/RegBank[11][15] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[11][13]  ( .G(n13142), .D(n13214), .Q(\pipeline/RegFile_DEC_WB/RegBank[11][13] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[11][0]  ( .G(n17716), .D(n13175), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[11][0] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[11][8]  ( .G(n17716), .D(n13199), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[11][8] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[11][14]  ( .G(n13142), .D(n13217), .Q(\pipeline/RegFile_DEC_WB/RegBank[11][14] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[11][16]  ( .G(n17716), .D(n13223), .Q(\pipeline/RegFile_DEC_WB/RegBank[11][16] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[11][18]  ( .G(n17716), .D(n13229), .Q(\pipeline/RegFile_DEC_WB/RegBank[11][18] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[11][20]  ( .G(n13142), .D(n13235), .Q(\pipeline/RegFile_DEC_WB/RegBank[11][20] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[11][22]  ( .G(n13142), .D(n13241), .Q(\pipeline/RegFile_DEC_WB/RegBank[11][22] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[11][24]  ( .G(n13142), .D(n13247), .Q(\pipeline/RegFile_DEC_WB/RegBank[11][24] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[11][26]  ( .G(n13142), .D(n13253), .Q(\pipeline/RegFile_DEC_WB/RegBank[11][26] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[11][28]  ( .G(n13142), .D(n13259), .Q(\pipeline/RegFile_DEC_WB/RegBank[11][28] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[11][30]  ( .G(n17716), .D(n13265), .Q(\pipeline/RegFile_DEC_WB/RegBank[11][30] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[12][31]  ( .G(n13139), .D(n13268), .Q(\pipeline/RegFile_DEC_WB/RegBank[12][31] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[12][29]  ( .G(n17717), .D(n13262), .Q(\pipeline/RegFile_DEC_WB/RegBank[12][29] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[12][27]  ( .G(n13139), .D(n13256), .Q(\pipeline/RegFile_DEC_WB/RegBank[12][27] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[12][25]  ( .G(n17717), .D(n13250), .Q(\pipeline/RegFile_DEC_WB/RegBank[12][25] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[12][23]  ( .G(n17717), .D(n13244), .Q(\pipeline/RegFile_DEC_WB/RegBank[12][23] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[12][21]  ( .G(n13139), .D(n13238), .Q(\pipeline/RegFile_DEC_WB/RegBank[12][21] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[12][19]  ( .G(n17717), .D(n13232), .Q(\pipeline/RegFile_DEC_WB/RegBank[12][19] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[12][17]  ( .G(n13139), .D(n13226), .Q(\pipeline/RegFile_DEC_WB/RegBank[12][17] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[12][15]  ( .G(n17717), .D(n13220), .Q(\pipeline/RegFile_DEC_WB/RegBank[12][15] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[12][13]  ( .G(n13139), .D(n13214), .Q(\pipeline/RegFile_DEC_WB/RegBank[12][13] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[12][0]  ( .G(n17717), .D(n13175), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[12][0] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[12][8]  ( .G(n17717), .D(n13199), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[12][8] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[12][14]  ( .G(n13139), .D(n13217), .Q(\pipeline/RegFile_DEC_WB/RegBank[12][14] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[12][16]  ( .G(n17717), .D(n13223), .Q(\pipeline/RegFile_DEC_WB/RegBank[12][16] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[12][18]  ( .G(n17717), .D(n13229), .Q(\pipeline/RegFile_DEC_WB/RegBank[12][18] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[12][20]  ( .G(n13139), .D(n13235), .Q(\pipeline/RegFile_DEC_WB/RegBank[12][20] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[12][22]  ( .G(n13139), .D(n13241), .Q(\pipeline/RegFile_DEC_WB/RegBank[12][22] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[12][24]  ( .G(n13139), .D(n13247), .Q(\pipeline/RegFile_DEC_WB/RegBank[12][24] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[12][26]  ( .G(n13139), .D(n13253), .Q(\pipeline/RegFile_DEC_WB/RegBank[12][26] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[12][28]  ( .G(n13139), .D(n13259), .Q(\pipeline/RegFile_DEC_WB/RegBank[12][28] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[12][30]  ( .G(n17717), .D(n13265), .Q(\pipeline/RegFile_DEC_WB/RegBank[12][30] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[13][31]  ( .G(n13136), .D(n13268), .Q(\pipeline/RegFile_DEC_WB/RegBank[13][31] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[13][29]  ( .G(n17718), .D(n13262), .Q(\pipeline/RegFile_DEC_WB/RegBank[13][29] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[13][27]  ( .G(n13136), .D(n13256), .Q(\pipeline/RegFile_DEC_WB/RegBank[13][27] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[13][25]  ( .G(n17718), .D(n13250), .Q(\pipeline/RegFile_DEC_WB/RegBank[13][25] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[13][23]  ( .G(n17718), .D(n13244), .Q(\pipeline/RegFile_DEC_WB/RegBank[13][23] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[13][21]  ( .G(n13136), .D(n13238), .Q(\pipeline/RegFile_DEC_WB/RegBank[13][21] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[13][19]  ( .G(n17718), .D(n13232), .Q(\pipeline/RegFile_DEC_WB/RegBank[13][19] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[13][17]  ( .G(n13136), .D(n13226), .Q(\pipeline/RegFile_DEC_WB/RegBank[13][17] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[13][15]  ( .G(n17718), .D(n13220), .Q(\pipeline/RegFile_DEC_WB/RegBank[13][15] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[13][13]  ( .G(n13136), .D(n13214), .Q(\pipeline/RegFile_DEC_WB/RegBank[13][13] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[13][0]  ( .G(n17718), .D(n13175), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[13][0] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[13][8]  ( .G(n17718), .D(n13199), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[13][8] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[13][14]  ( .G(n13136), .D(n13217), .Q(\pipeline/RegFile_DEC_WB/RegBank[13][14] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[13][16]  ( .G(n17718), .D(n13223), .Q(\pipeline/RegFile_DEC_WB/RegBank[13][16] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[13][18]  ( .G(n17718), .D(n13229), .Q(\pipeline/RegFile_DEC_WB/RegBank[13][18] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[13][20]  ( .G(n13136), .D(n13235), .Q(\pipeline/RegFile_DEC_WB/RegBank[13][20] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[13][22]  ( .G(n13136), .D(n13241), .Q(\pipeline/RegFile_DEC_WB/RegBank[13][22] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[13][24]  ( .G(n13136), .D(n13247), .Q(\pipeline/RegFile_DEC_WB/RegBank[13][24] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[13][26]  ( .G(n13136), .D(n13253), .Q(\pipeline/RegFile_DEC_WB/RegBank[13][26] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[13][28]  ( .G(n13136), .D(n13259), .Q(\pipeline/RegFile_DEC_WB/RegBank[13][28] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[13][30]  ( .G(n17718), .D(n13265), .Q(\pipeline/RegFile_DEC_WB/RegBank[13][30] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[14][31]  ( .G(n13133), .D(n13268), .Q(\pipeline/RegFile_DEC_WB/RegBank[14][31] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[14][29]  ( .G(n17719), .D(n13262), .Q(\pipeline/RegFile_DEC_WB/RegBank[14][29] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[14][27]  ( .G(n13133), .D(n13256), .Q(\pipeline/RegFile_DEC_WB/RegBank[14][27] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[14][25]  ( .G(n17719), .D(n13250), .Q(\pipeline/RegFile_DEC_WB/RegBank[14][25] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[14][23]  ( .G(n17719), .D(n13244), .Q(\pipeline/RegFile_DEC_WB/RegBank[14][23] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[14][21]  ( .G(n13133), .D(n13238), .Q(\pipeline/RegFile_DEC_WB/RegBank[14][21] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[14][19]  ( .G(n17719), .D(n13232), .Q(\pipeline/RegFile_DEC_WB/RegBank[14][19] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[14][17]  ( .G(n13133), .D(n13226), .Q(\pipeline/RegFile_DEC_WB/RegBank[14][17] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[14][15]  ( .G(n17719), .D(n13220), .Q(\pipeline/RegFile_DEC_WB/RegBank[14][15] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[14][13]  ( .G(n13133), .D(n13214), .Q(\pipeline/RegFile_DEC_WB/RegBank[14][13] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[14][0]  ( .G(n17719), .D(n13175), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[14][0] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[14][8]  ( .G(n17719), .D(n13199), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[14][8] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[14][14]  ( .G(n13133), .D(n13217), .Q(\pipeline/RegFile_DEC_WB/RegBank[14][14] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[14][16]  ( .G(n17719), .D(n13223), .Q(\pipeline/RegFile_DEC_WB/RegBank[14][16] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[14][18]  ( .G(n17719), .D(n13229), .Q(\pipeline/RegFile_DEC_WB/RegBank[14][18] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[14][20]  ( .G(n13133), .D(n13235), .Q(\pipeline/RegFile_DEC_WB/RegBank[14][20] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[14][22]  ( .G(n13133), .D(n13241), .Q(\pipeline/RegFile_DEC_WB/RegBank[14][22] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[14][24]  ( .G(n13133), .D(n13247), .Q(\pipeline/RegFile_DEC_WB/RegBank[14][24] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[14][26]  ( .G(n13133), .D(n13253), .Q(\pipeline/RegFile_DEC_WB/RegBank[14][26] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[14][28]  ( .G(n13133), .D(n13259), .Q(\pipeline/RegFile_DEC_WB/RegBank[14][28] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[14][30]  ( .G(n17719), .D(n13265), .Q(\pipeline/RegFile_DEC_WB/RegBank[14][30] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[15][31]  ( .G(n13130), .D(n13268), .Q(\pipeline/RegFile_DEC_WB/RegBank[15][31] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[15][29]  ( .G(n17720), .D(n13262), .Q(\pipeline/RegFile_DEC_WB/RegBank[15][29] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[15][27]  ( .G(n13130), .D(n13256), .Q(\pipeline/RegFile_DEC_WB/RegBank[15][27] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[15][25]  ( .G(n17720), .D(n13250), .Q(\pipeline/RegFile_DEC_WB/RegBank[15][25] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[15][23]  ( .G(n17720), .D(n13244), .Q(\pipeline/RegFile_DEC_WB/RegBank[15][23] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[15][21]  ( .G(n13130), .D(n13238), .Q(\pipeline/RegFile_DEC_WB/RegBank[15][21] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[15][19]  ( .G(n17720), .D(n13232), .Q(\pipeline/RegFile_DEC_WB/RegBank[15][19] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[15][17]  ( .G(n13130), .D(n13226), .Q(\pipeline/RegFile_DEC_WB/RegBank[15][17] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[15][15]  ( .G(n17720), .D(n13220), .Q(\pipeline/RegFile_DEC_WB/RegBank[15][15] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[15][13]  ( .G(n13130), .D(n13214), .Q(\pipeline/RegFile_DEC_WB/RegBank[15][13] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[15][0]  ( .G(n17720), .D(n13175), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[15][0] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[15][8]  ( .G(n17720), .D(n13199), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[15][8] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[15][14]  ( .G(n13130), .D(n13217), .Q(\pipeline/RegFile_DEC_WB/RegBank[15][14] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[15][16]  ( .G(n17720), .D(n13223), .Q(\pipeline/RegFile_DEC_WB/RegBank[15][16] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[15][18]  ( .G(n17720), .D(n13229), .Q(\pipeline/RegFile_DEC_WB/RegBank[15][18] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[15][20]  ( .G(n13130), .D(n13235), .Q(\pipeline/RegFile_DEC_WB/RegBank[15][20] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[15][22]  ( .G(n13130), .D(n13241), .Q(\pipeline/RegFile_DEC_WB/RegBank[15][22] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[15][24]  ( .G(n13130), .D(n13247), .Q(\pipeline/RegFile_DEC_WB/RegBank[15][24] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[15][26]  ( .G(n13130), .D(n13253), .Q(\pipeline/RegFile_DEC_WB/RegBank[15][26] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[15][28]  ( .G(n13130), .D(n13259), .Q(\pipeline/RegFile_DEC_WB/RegBank[15][28] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[15][30]  ( .G(n17720), .D(n13265), .Q(\pipeline/RegFile_DEC_WB/RegBank[15][30] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[16][31]  ( .G(n13127), .D(n13268), .Q(\pipeline/RegFile_DEC_WB/RegBank[16][31] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[16][29]  ( .G(n17721), .D(n13262), .Q(\pipeline/RegFile_DEC_WB/RegBank[16][29] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[16][27]  ( .G(n13127), .D(n13256), .Q(\pipeline/RegFile_DEC_WB/RegBank[16][27] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[16][25]  ( .G(n17721), .D(n13250), .Q(\pipeline/RegFile_DEC_WB/RegBank[16][25] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[16][23]  ( .G(n17721), .D(n13244), .Q(\pipeline/RegFile_DEC_WB/RegBank[16][23] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[16][21]  ( .G(n13127), .D(n13238), .Q(\pipeline/RegFile_DEC_WB/RegBank[16][21] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[16][19]  ( .G(n17721), .D(n13232), .Q(\pipeline/RegFile_DEC_WB/RegBank[16][19] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[16][17]  ( .G(n13127), .D(n13226), .Q(\pipeline/RegFile_DEC_WB/RegBank[16][17] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[16][15]  ( .G(n17721), .D(n13220), .Q(\pipeline/RegFile_DEC_WB/RegBank[16][15] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[16][13]  ( .G(n13127), .D(n13214), .Q(\pipeline/RegFile_DEC_WB/RegBank[16][13] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[16][0]  ( .G(n17721), .D(n13175), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[16][0] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[16][8]  ( .G(n17721), .D(n13199), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[16][8] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[16][14]  ( .G(n13127), .D(n13217), .Q(\pipeline/RegFile_DEC_WB/RegBank[16][14] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[16][16]  ( .G(n17721), .D(n13223), .Q(\pipeline/RegFile_DEC_WB/RegBank[16][16] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[16][18]  ( .G(n17721), .D(n13229), .Q(\pipeline/RegFile_DEC_WB/RegBank[16][18] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[16][20]  ( .G(n13127), .D(n13235), .Q(\pipeline/RegFile_DEC_WB/RegBank[16][20] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[16][22]  ( .G(n13127), .D(n13241), .Q(\pipeline/RegFile_DEC_WB/RegBank[16][22] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[16][24]  ( .G(n13127), .D(n13247), .Q(\pipeline/RegFile_DEC_WB/RegBank[16][24] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[16][26]  ( .G(n13127), .D(n13253), .Q(\pipeline/RegFile_DEC_WB/RegBank[16][26] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[16][28]  ( .G(n13127), .D(n13259), .Q(\pipeline/RegFile_DEC_WB/RegBank[16][28] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[16][30]  ( .G(n17721), .D(n13265), .Q(\pipeline/RegFile_DEC_WB/RegBank[16][30] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[17][31]  ( .G(n13124), .D(n13268), .Q(\pipeline/RegFile_DEC_WB/RegBank[17][31] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[17][29]  ( .G(n17722), .D(n13262), .Q(\pipeline/RegFile_DEC_WB/RegBank[17][29] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[17][27]  ( .G(n13124), .D(n13256), .Q(\pipeline/RegFile_DEC_WB/RegBank[17][27] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[17][25]  ( .G(n17722), .D(n13250), .Q(\pipeline/RegFile_DEC_WB/RegBank[17][25] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[17][23]  ( .G(n17722), .D(n13244), .Q(\pipeline/RegFile_DEC_WB/RegBank[17][23] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[17][21]  ( .G(n13124), .D(n13238), .Q(\pipeline/RegFile_DEC_WB/RegBank[17][21] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[17][19]  ( .G(n17722), .D(n13232), .Q(\pipeline/RegFile_DEC_WB/RegBank[17][19] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[17][17]  ( .G(n13124), .D(n13226), .Q(\pipeline/RegFile_DEC_WB/RegBank[17][17] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[17][15]  ( .G(n17722), .D(n13220), .Q(\pipeline/RegFile_DEC_WB/RegBank[17][15] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[17][13]  ( .G(n13124), .D(n13214), .Q(\pipeline/RegFile_DEC_WB/RegBank[17][13] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[17][0]  ( .G(n17722), .D(n13175), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[17][0] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[17][8]  ( .G(n17722), .D(n13199), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[17][8] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[17][14]  ( .G(n13124), .D(n13217), .Q(\pipeline/RegFile_DEC_WB/RegBank[17][14] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[17][16]  ( .G(n17722), .D(n13223), .Q(\pipeline/RegFile_DEC_WB/RegBank[17][16] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[17][18]  ( .G(n17722), .D(n13229), .Q(\pipeline/RegFile_DEC_WB/RegBank[17][18] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[17][20]  ( .G(n13124), .D(n13235), .Q(\pipeline/RegFile_DEC_WB/RegBank[17][20] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[17][22]  ( .G(n13124), .D(n13241), .Q(\pipeline/RegFile_DEC_WB/RegBank[17][22] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[17][24]  ( .G(n13124), .D(n13247), .Q(\pipeline/RegFile_DEC_WB/RegBank[17][24] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[17][26]  ( .G(n13124), .D(n13253), .Q(\pipeline/RegFile_DEC_WB/RegBank[17][26] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[17][28]  ( .G(n13124), .D(n13259), .Q(\pipeline/RegFile_DEC_WB/RegBank[17][28] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[17][30]  ( .G(n17722), .D(n13265), .Q(\pipeline/RegFile_DEC_WB/RegBank[17][30] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[18][31]  ( .G(n13121), .D(n13268), .Q(\pipeline/RegFile_DEC_WB/RegBank[18][31] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[18][29]  ( .G(n17723), .D(n13262), .Q(\pipeline/RegFile_DEC_WB/RegBank[18][29] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[18][27]  ( .G(n13121), .D(n13256), .Q(\pipeline/RegFile_DEC_WB/RegBank[18][27] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[18][25]  ( .G(n17723), .D(n13250), .Q(\pipeline/RegFile_DEC_WB/RegBank[18][25] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[18][23]  ( .G(n17723), .D(n13244), .Q(\pipeline/RegFile_DEC_WB/RegBank[18][23] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[18][21]  ( .G(n13121), .D(n13238), .Q(\pipeline/RegFile_DEC_WB/RegBank[18][21] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[18][19]  ( .G(n17723), .D(n13232), .Q(\pipeline/RegFile_DEC_WB/RegBank[18][19] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[18][17]  ( .G(n13121), .D(n13226), .Q(\pipeline/RegFile_DEC_WB/RegBank[18][17] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[18][15]  ( .G(n17723), .D(n13220), .Q(\pipeline/RegFile_DEC_WB/RegBank[18][15] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[18][13]  ( .G(n13121), .D(n13214), .Q(\pipeline/RegFile_DEC_WB/RegBank[18][13] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[18][0]  ( .G(n17723), .D(n13175), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[18][0] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[18][8]  ( .G(n17723), .D(n13199), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[18][8] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[18][14]  ( .G(n13121), .D(n13217), .Q(\pipeline/RegFile_DEC_WB/RegBank[18][14] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[18][16]  ( .G(n17723), .D(n13223), .Q(\pipeline/RegFile_DEC_WB/RegBank[18][16] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[18][18]  ( .G(n17723), .D(n13229), .Q(\pipeline/RegFile_DEC_WB/RegBank[18][18] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[18][20]  ( .G(n13121), .D(n13235), .Q(\pipeline/RegFile_DEC_WB/RegBank[18][20] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[18][22]  ( .G(n13121), .D(n13241), .Q(\pipeline/RegFile_DEC_WB/RegBank[18][22] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[18][24]  ( .G(n13121), .D(n13247), .Q(\pipeline/RegFile_DEC_WB/RegBank[18][24] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[18][26]  ( .G(n13121), .D(n13253), .Q(\pipeline/RegFile_DEC_WB/RegBank[18][26] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[18][28]  ( .G(n13121), .D(n13259), .Q(\pipeline/RegFile_DEC_WB/RegBank[18][28] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[18][30]  ( .G(n17723), .D(n13265), .Q(\pipeline/RegFile_DEC_WB/RegBank[18][30] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[19][31]  ( .G(n13118), .D(n13268), .Q(\pipeline/RegFile_DEC_WB/RegBank[19][31] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[19][29]  ( .G(n17724), .D(n13262), .Q(\pipeline/RegFile_DEC_WB/RegBank[19][29] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[19][27]  ( .G(n13118), .D(n13256), .Q(\pipeline/RegFile_DEC_WB/RegBank[19][27] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[19][25]  ( .G(n17724), .D(n13250), .Q(\pipeline/RegFile_DEC_WB/RegBank[19][25] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[19][23]  ( .G(n17724), .D(n13244), .Q(\pipeline/RegFile_DEC_WB/RegBank[19][23] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[19][21]  ( .G(n13118), .D(n13238), .Q(\pipeline/RegFile_DEC_WB/RegBank[19][21] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[19][19]  ( .G(n17724), .D(n13232), .Q(\pipeline/RegFile_DEC_WB/RegBank[19][19] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[19][17]  ( .G(n13118), .D(n13226), .Q(\pipeline/RegFile_DEC_WB/RegBank[19][17] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[19][15]  ( .G(n17724), .D(n13220), .Q(\pipeline/RegFile_DEC_WB/RegBank[19][15] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[19][13]  ( .G(n13118), .D(n13214), .Q(\pipeline/RegFile_DEC_WB/RegBank[19][13] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[19][0]  ( .G(n17724), .D(n13175), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[19][0] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[19][8]  ( .G(n17724), .D(n13199), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[19][8] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[19][14]  ( .G(n13118), .D(n13217), .Q(\pipeline/RegFile_DEC_WB/RegBank[19][14] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[19][16]  ( .G(n17724), .D(n13223), .Q(\pipeline/RegFile_DEC_WB/RegBank[19][16] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[19][18]  ( .G(n17724), .D(n13229), .Q(\pipeline/RegFile_DEC_WB/RegBank[19][18] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[19][20]  ( .G(n13118), .D(n13235), .Q(\pipeline/RegFile_DEC_WB/RegBank[19][20] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[19][22]  ( .G(n13118), .D(n13241), .Q(\pipeline/RegFile_DEC_WB/RegBank[19][22] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[19][24]  ( .G(n13118), .D(n13247), .Q(\pipeline/RegFile_DEC_WB/RegBank[19][24] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[19][26]  ( .G(n13118), .D(n13253), .Q(\pipeline/RegFile_DEC_WB/RegBank[19][26] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[19][28]  ( .G(n13118), .D(n13259), .Q(\pipeline/RegFile_DEC_WB/RegBank[19][28] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[19][30]  ( .G(n17724), .D(n13265), .Q(\pipeline/RegFile_DEC_WB/RegBank[19][30] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[20][31]  ( .G(n13115), .D(n13268), .Q(\pipeline/RegFile_DEC_WB/RegBank[20][31] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[20][29]  ( .G(n17725), .D(n13262), .Q(\pipeline/RegFile_DEC_WB/RegBank[20][29] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[20][27]  ( .G(n13115), .D(n13256), .Q(\pipeline/RegFile_DEC_WB/RegBank[20][27] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[20][25]  ( .G(n17725), .D(n13250), .Q(\pipeline/RegFile_DEC_WB/RegBank[20][25] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[20][23]  ( .G(n17725), .D(n13244), .Q(\pipeline/RegFile_DEC_WB/RegBank[20][23] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[20][21]  ( .G(n13115), .D(n13238), .Q(\pipeline/RegFile_DEC_WB/RegBank[20][21] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[20][19]  ( .G(n17725), .D(n13232), .Q(\pipeline/RegFile_DEC_WB/RegBank[20][19] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[20][17]  ( .G(n13115), .D(n13226), .Q(\pipeline/RegFile_DEC_WB/RegBank[20][17] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[20][15]  ( .G(n17725), .D(n13220), .Q(\pipeline/RegFile_DEC_WB/RegBank[20][15] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[20][13]  ( .G(n13115), .D(n13214), .Q(\pipeline/RegFile_DEC_WB/RegBank[20][13] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[20][0]  ( .G(n17725), .D(n13175), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[20][0] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[20][8]  ( .G(n17725), .D(n13199), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[20][8] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[20][14]  ( .G(n13115), .D(n13217), .Q(\pipeline/RegFile_DEC_WB/RegBank[20][14] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[20][16]  ( .G(n17725), .D(n13223), .Q(\pipeline/RegFile_DEC_WB/RegBank[20][16] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[20][18]  ( .G(n17725), .D(n13229), .Q(\pipeline/RegFile_DEC_WB/RegBank[20][18] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[20][20]  ( .G(n13115), .D(n13235), .Q(\pipeline/RegFile_DEC_WB/RegBank[20][20] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[20][22]  ( .G(n13115), .D(n13241), .Q(\pipeline/RegFile_DEC_WB/RegBank[20][22] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[20][24]  ( .G(n13115), .D(n13247), .Q(\pipeline/RegFile_DEC_WB/RegBank[20][24] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[20][26]  ( .G(n13115), .D(n13253), .Q(\pipeline/RegFile_DEC_WB/RegBank[20][26] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[20][28]  ( .G(n13115), .D(n13259), .Q(\pipeline/RegFile_DEC_WB/RegBank[20][28] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[20][30]  ( .G(n17725), .D(n13265), .Q(\pipeline/RegFile_DEC_WB/RegBank[20][30] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[21][31]  ( .G(n13112), .D(n13268), .Q(\pipeline/RegFile_DEC_WB/RegBank[21][31] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[21][29]  ( .G(n17726), .D(n13262), .Q(\pipeline/RegFile_DEC_WB/RegBank[21][29] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[21][27]  ( .G(n13112), .D(n13256), .Q(\pipeline/RegFile_DEC_WB/RegBank[21][27] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[21][25]  ( .G(n17726), .D(n13250), .Q(\pipeline/RegFile_DEC_WB/RegBank[21][25] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[21][23]  ( .G(n17726), .D(n13244), .Q(\pipeline/RegFile_DEC_WB/RegBank[21][23] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[21][21]  ( .G(n13112), .D(n13238), .Q(\pipeline/RegFile_DEC_WB/RegBank[21][21] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[21][19]  ( .G(n17726), .D(n13232), .Q(\pipeline/RegFile_DEC_WB/RegBank[21][19] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[21][17]  ( .G(n13112), .D(n13226), .Q(\pipeline/RegFile_DEC_WB/RegBank[21][17] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[21][15]  ( .G(n17726), .D(n13220), .Q(\pipeline/RegFile_DEC_WB/RegBank[21][15] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[21][13]  ( .G(n13112), .D(n13214), .Q(\pipeline/RegFile_DEC_WB/RegBank[21][13] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[21][0]  ( .G(n17726), .D(n13175), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[21][0] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[21][8]  ( .G(n17726), .D(n13199), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[21][8] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[21][14]  ( .G(n13112), .D(n13217), .Q(\pipeline/RegFile_DEC_WB/RegBank[21][14] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[21][16]  ( .G(n17726), .D(n13223), .Q(\pipeline/RegFile_DEC_WB/RegBank[21][16] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[21][18]  ( .G(n17726), .D(n13229), .Q(\pipeline/RegFile_DEC_WB/RegBank[21][18] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[21][20]  ( .G(n13112), .D(n13235), .Q(\pipeline/RegFile_DEC_WB/RegBank[21][20] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[21][22]  ( .G(n13112), .D(n13241), .Q(\pipeline/RegFile_DEC_WB/RegBank[21][22] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[21][24]  ( .G(n13112), .D(n13247), .Q(\pipeline/RegFile_DEC_WB/RegBank[21][24] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[21][26]  ( .G(n13112), .D(n13253), .Q(\pipeline/RegFile_DEC_WB/RegBank[21][26] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[21][28]  ( .G(n13112), .D(n13259), .Q(\pipeline/RegFile_DEC_WB/RegBank[21][28] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[21][30]  ( .G(n17726), .D(n13265), .Q(\pipeline/RegFile_DEC_WB/RegBank[21][30] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[22][31]  ( .G(n13109), .D(n13268), .Q(\pipeline/RegFile_DEC_WB/RegBank[22][31] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[22][29]  ( .G(n17727), .D(n13262), .Q(\pipeline/RegFile_DEC_WB/RegBank[22][29] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[22][27]  ( .G(n13109), .D(n13256), .Q(\pipeline/RegFile_DEC_WB/RegBank[22][27] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[22][25]  ( .G(n17727), .D(n13250), .Q(\pipeline/RegFile_DEC_WB/RegBank[22][25] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[22][23]  ( .G(n17727), .D(n13244), .Q(\pipeline/RegFile_DEC_WB/RegBank[22][23] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[22][21]  ( .G(n13109), .D(n13238), .Q(\pipeline/RegFile_DEC_WB/RegBank[22][21] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[22][19]  ( .G(n17727), .D(n13232), .Q(\pipeline/RegFile_DEC_WB/RegBank[22][19] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[22][17]  ( .G(n13109), .D(n13226), .Q(\pipeline/RegFile_DEC_WB/RegBank[22][17] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[22][15]  ( .G(n17727), .D(n13220), .Q(\pipeline/RegFile_DEC_WB/RegBank[22][15] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[22][13]  ( .G(n13109), .D(n13214), .Q(\pipeline/RegFile_DEC_WB/RegBank[22][13] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[22][0]  ( .G(n17727), .D(n13175), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[22][0] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[22][8]  ( .G(n17727), .D(n13199), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[22][8] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[22][14]  ( .G(n13109), .D(n13217), .Q(\pipeline/RegFile_DEC_WB/RegBank[22][14] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[22][16]  ( .G(n17727), .D(n13223), .Q(\pipeline/RegFile_DEC_WB/RegBank[22][16] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[22][18]  ( .G(n17727), .D(n13229), .Q(\pipeline/RegFile_DEC_WB/RegBank[22][18] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[22][20]  ( .G(n13109), .D(n13235), .Q(\pipeline/RegFile_DEC_WB/RegBank[22][20] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[22][22]  ( .G(n13109), .D(n13241), .Q(\pipeline/RegFile_DEC_WB/RegBank[22][22] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[22][24]  ( .G(n13109), .D(n13247), .Q(\pipeline/RegFile_DEC_WB/RegBank[22][24] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[22][26]  ( .G(n13109), .D(n13253), .Q(\pipeline/RegFile_DEC_WB/RegBank[22][26] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[22][28]  ( .G(n13109), .D(n13259), .Q(\pipeline/RegFile_DEC_WB/RegBank[22][28] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[22][30]  ( .G(n17727), .D(n13265), .Q(\pipeline/RegFile_DEC_WB/RegBank[22][30] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[23][31]  ( .G(n13106), .D(n13268), .Q(\pipeline/RegFile_DEC_WB/RegBank[23][31] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[23][29]  ( .G(n17728), .D(n13262), .Q(\pipeline/RegFile_DEC_WB/RegBank[23][29] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[23][27]  ( .G(n13106), .D(n13256), .Q(\pipeline/RegFile_DEC_WB/RegBank[23][27] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[23][25]  ( .G(n17728), .D(n13250), .Q(\pipeline/RegFile_DEC_WB/RegBank[23][25] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[23][23]  ( .G(n17728), .D(n13244), .Q(\pipeline/RegFile_DEC_WB/RegBank[23][23] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[23][21]  ( .G(n13106), .D(n13238), .Q(\pipeline/RegFile_DEC_WB/RegBank[23][21] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[23][19]  ( .G(n17728), .D(n13232), .Q(\pipeline/RegFile_DEC_WB/RegBank[23][19] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[23][17]  ( .G(n13106), .D(n13226), .Q(\pipeline/RegFile_DEC_WB/RegBank[23][17] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[23][15]  ( .G(n17728), .D(n13220), .Q(\pipeline/RegFile_DEC_WB/RegBank[23][15] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[23][13]  ( .G(n13106), .D(n13214), .Q(\pipeline/RegFile_DEC_WB/RegBank[23][13] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[23][0]  ( .G(n17728), .D(n13175), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[23][0] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[23][8]  ( .G(n17728), .D(n13199), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[23][8] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[23][14]  ( .G(n13106), .D(n13217), .Q(\pipeline/RegFile_DEC_WB/RegBank[23][14] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[23][16]  ( .G(n17728), .D(n13223), .Q(\pipeline/RegFile_DEC_WB/RegBank[23][16] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[23][18]  ( .G(n17728), .D(n13229), .Q(\pipeline/RegFile_DEC_WB/RegBank[23][18] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[23][20]  ( .G(n13106), .D(n13235), .Q(\pipeline/RegFile_DEC_WB/RegBank[23][20] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[23][22]  ( .G(n13106), .D(n13241), .Q(\pipeline/RegFile_DEC_WB/RegBank[23][22] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[23][24]  ( .G(n13106), .D(n13247), .Q(\pipeline/RegFile_DEC_WB/RegBank[23][24] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[23][26]  ( .G(n13106), .D(n13253), .Q(\pipeline/RegFile_DEC_WB/RegBank[23][26] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[23][28]  ( .G(n13106), .D(n13259), .Q(\pipeline/RegFile_DEC_WB/RegBank[23][28] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[23][30]  ( .G(n17728), .D(n13265), .Q(\pipeline/RegFile_DEC_WB/RegBank[23][30] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[24][31]  ( .G(n13103), .D(n13268), .Q(\pipeline/RegFile_DEC_WB/RegBank[24][31] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[24][29]  ( .G(n17729), .D(n13262), .Q(\pipeline/RegFile_DEC_WB/RegBank[24][29] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[24][27]  ( .G(n13103), .D(n13256), .Q(\pipeline/RegFile_DEC_WB/RegBank[24][27] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[24][25]  ( .G(n17729), .D(n13250), .Q(\pipeline/RegFile_DEC_WB/RegBank[24][25] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[24][23]  ( .G(n17729), .D(n13244), .Q(\pipeline/RegFile_DEC_WB/RegBank[24][23] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[24][21]  ( .G(n13103), .D(n13238), .Q(\pipeline/RegFile_DEC_WB/RegBank[24][21] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[24][19]  ( .G(n17729), .D(n13232), .Q(\pipeline/RegFile_DEC_WB/RegBank[24][19] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[24][17]  ( .G(n13103), .D(n13226), .Q(\pipeline/RegFile_DEC_WB/RegBank[24][17] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[24][15]  ( .G(n17729), .D(n13220), .Q(\pipeline/RegFile_DEC_WB/RegBank[24][15] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[24][13]  ( .G(n13103), .D(n13214), .Q(\pipeline/RegFile_DEC_WB/RegBank[24][13] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[24][0]  ( .G(n17729), .D(n13175), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[24][0] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[24][8]  ( .G(n17729), .D(n13199), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[24][8] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[24][14]  ( .G(n13103), .D(n13217), .Q(\pipeline/RegFile_DEC_WB/RegBank[24][14] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[24][16]  ( .G(n17729), .D(n13223), .Q(\pipeline/RegFile_DEC_WB/RegBank[24][16] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[24][18]  ( .G(n17729), .D(n13229), .Q(\pipeline/RegFile_DEC_WB/RegBank[24][18] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[24][20]  ( .G(n13103), .D(n13235), .Q(\pipeline/RegFile_DEC_WB/RegBank[24][20] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[24][22]  ( .G(n13103), .D(n13241), .Q(\pipeline/RegFile_DEC_WB/RegBank[24][22] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[24][24]  ( .G(n13103), .D(n13247), .Q(\pipeline/RegFile_DEC_WB/RegBank[24][24] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[24][26]  ( .G(n13103), .D(n13253), .Q(\pipeline/RegFile_DEC_WB/RegBank[24][26] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[24][28]  ( .G(n13103), .D(n13259), .Q(\pipeline/RegFile_DEC_WB/RegBank[24][28] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[24][30]  ( .G(n17729), .D(n13265), .Q(\pipeline/RegFile_DEC_WB/RegBank[24][30] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[25][31]  ( .G(n13100), .D(n13268), .Q(\pipeline/RegFile_DEC_WB/RegBank[25][31] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[25][29]  ( .G(n17730), .D(n13262), .Q(\pipeline/RegFile_DEC_WB/RegBank[25][29] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[25][27]  ( .G(n13100), .D(n13256), .Q(\pipeline/RegFile_DEC_WB/RegBank[25][27] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[25][25]  ( .G(n17730), .D(n13250), .Q(\pipeline/RegFile_DEC_WB/RegBank[25][25] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[25][23]  ( .G(n17730), .D(n13244), .Q(\pipeline/RegFile_DEC_WB/RegBank[25][23] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[25][21]  ( .G(n13100), .D(n13238), .Q(\pipeline/RegFile_DEC_WB/RegBank[25][21] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[25][19]  ( .G(n17730), .D(n13232), .Q(\pipeline/RegFile_DEC_WB/RegBank[25][19] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[25][17]  ( .G(n13100), .D(n13226), .Q(\pipeline/RegFile_DEC_WB/RegBank[25][17] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[25][15]  ( .G(n17730), .D(n13220), .Q(\pipeline/RegFile_DEC_WB/RegBank[25][15] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[25][13]  ( .G(n13100), .D(n13214), .Q(\pipeline/RegFile_DEC_WB/RegBank[25][13] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[25][0]  ( .G(n17730), .D(n13175), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[25][0] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[25][8]  ( .G(n17730), .D(n13199), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[25][8] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[25][14]  ( .G(n13100), .D(n13217), .Q(\pipeline/RegFile_DEC_WB/RegBank[25][14] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[25][16]  ( .G(n17730), .D(n13223), .Q(\pipeline/RegFile_DEC_WB/RegBank[25][16] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[25][18]  ( .G(n17730), .D(n13229), .Q(\pipeline/RegFile_DEC_WB/RegBank[25][18] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[25][20]  ( .G(n13100), .D(n13235), .Q(\pipeline/RegFile_DEC_WB/RegBank[25][20] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[25][22]  ( .G(n13100), .D(n13241), .Q(\pipeline/RegFile_DEC_WB/RegBank[25][22] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[25][24]  ( .G(n13100), .D(n13247), .Q(\pipeline/RegFile_DEC_WB/RegBank[25][24] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[25][26]  ( .G(n13100), .D(n13253), .Q(\pipeline/RegFile_DEC_WB/RegBank[25][26] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[25][28]  ( .G(n13100), .D(n13259), .Q(\pipeline/RegFile_DEC_WB/RegBank[25][28] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[25][30]  ( .G(n17730), .D(n13265), .Q(\pipeline/RegFile_DEC_WB/RegBank[25][30] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[26][31]  ( .G(n13097), .D(n13268), .Q(\pipeline/RegFile_DEC_WB/RegBank[26][31] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[26][29]  ( .G(n17731), .D(n13262), .Q(\pipeline/RegFile_DEC_WB/RegBank[26][29] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[26][27]  ( .G(n13097), .D(n13256), .Q(\pipeline/RegFile_DEC_WB/RegBank[26][27] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[26][25]  ( .G(n17731), .D(n13250), .Q(\pipeline/RegFile_DEC_WB/RegBank[26][25] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[26][23]  ( .G(n17731), .D(n13244), .Q(\pipeline/RegFile_DEC_WB/RegBank[26][23] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[26][21]  ( .G(n13097), .D(n13238), .Q(\pipeline/RegFile_DEC_WB/RegBank[26][21] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[26][19]  ( .G(n17731), .D(n13232), .Q(\pipeline/RegFile_DEC_WB/RegBank[26][19] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[26][17]  ( .G(n13097), .D(n13226), .Q(\pipeline/RegFile_DEC_WB/RegBank[26][17] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[26][15]  ( .G(n17731), .D(n13220), .Q(\pipeline/RegFile_DEC_WB/RegBank[26][15] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[26][13]  ( .G(n13097), .D(n13214), .Q(\pipeline/RegFile_DEC_WB/RegBank[26][13] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[26][0]  ( .G(n17731), .D(n13175), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[26][0] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[26][8]  ( .G(n17731), .D(n13199), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[26][8] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[26][14]  ( .G(n13097), .D(n13217), .Q(\pipeline/RegFile_DEC_WB/RegBank[26][14] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[26][16]  ( .G(n17731), .D(n13223), .Q(\pipeline/RegFile_DEC_WB/RegBank[26][16] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[26][18]  ( .G(n17731), .D(n13229), .Q(\pipeline/RegFile_DEC_WB/RegBank[26][18] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[26][20]  ( .G(n13097), .D(n13235), .Q(\pipeline/RegFile_DEC_WB/RegBank[26][20] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[26][22]  ( .G(n13097), .D(n13241), .Q(\pipeline/RegFile_DEC_WB/RegBank[26][22] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[26][24]  ( .G(n13097), .D(n13247), .Q(\pipeline/RegFile_DEC_WB/RegBank[26][24] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[26][26]  ( .G(n13097), .D(n13253), .Q(\pipeline/RegFile_DEC_WB/RegBank[26][26] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[26][28]  ( .G(n13097), .D(n13259), .Q(\pipeline/RegFile_DEC_WB/RegBank[26][28] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[26][30]  ( .G(n17731), .D(n13265), .Q(\pipeline/RegFile_DEC_WB/RegBank[26][30] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[27][31]  ( .G(n13094), .D(n13268), .Q(\pipeline/RegFile_DEC_WB/RegBank[27][31] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[27][29]  ( .G(n17732), .D(n13262), .Q(\pipeline/RegFile_DEC_WB/RegBank[27][29] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[27][27]  ( .G(n13094), .D(n13256), .Q(\pipeline/RegFile_DEC_WB/RegBank[27][27] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[27][25]  ( .G(n17732), .D(n13250), .Q(\pipeline/RegFile_DEC_WB/RegBank[27][25] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[27][23]  ( .G(n17732), .D(n13244), .Q(\pipeline/RegFile_DEC_WB/RegBank[27][23] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[27][21]  ( .G(n13094), .D(n13238), .Q(\pipeline/RegFile_DEC_WB/RegBank[27][21] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[27][19]  ( .G(n17732), .D(n13232), .Q(\pipeline/RegFile_DEC_WB/RegBank[27][19] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[27][17]  ( .G(n13094), .D(n13226), .Q(\pipeline/RegFile_DEC_WB/RegBank[27][17] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[27][15]  ( .G(n17732), .D(n13220), .Q(\pipeline/RegFile_DEC_WB/RegBank[27][15] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[27][13]  ( .G(n13094), .D(n13214), .Q(\pipeline/RegFile_DEC_WB/RegBank[27][13] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[27][0]  ( .G(n17732), .D(n13175), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[27][0] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[27][8]  ( .G(n17732), .D(n13199), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[27][8] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[27][14]  ( .G(n13094), .D(n13217), .Q(\pipeline/RegFile_DEC_WB/RegBank[27][14] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[27][16]  ( .G(n17732), .D(n13223), .Q(\pipeline/RegFile_DEC_WB/RegBank[27][16] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[27][18]  ( .G(n17732), .D(n13229), .Q(\pipeline/RegFile_DEC_WB/RegBank[27][18] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[27][20]  ( .G(n13094), .D(n13235), .Q(\pipeline/RegFile_DEC_WB/RegBank[27][20] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[27][22]  ( .G(n13094), .D(n13241), .Q(\pipeline/RegFile_DEC_WB/RegBank[27][22] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[27][24]  ( .G(n13094), .D(n13247), .Q(\pipeline/RegFile_DEC_WB/RegBank[27][24] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[27][26]  ( .G(n13094), .D(n13253), .Q(\pipeline/RegFile_DEC_WB/RegBank[27][26] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[27][28]  ( .G(n13094), .D(n13259), .Q(\pipeline/RegFile_DEC_WB/RegBank[27][28] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[27][30]  ( .G(n17732), .D(n13265), .Q(\pipeline/RegFile_DEC_WB/RegBank[27][30] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[28][31]  ( .G(n13091), .D(n13268), .Q(\pipeline/RegFile_DEC_WB/RegBank[28][31] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[28][29]  ( .G(n17733), .D(n13262), .Q(\pipeline/RegFile_DEC_WB/RegBank[28][29] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[28][27]  ( .G(n13091), .D(n13256), .Q(\pipeline/RegFile_DEC_WB/RegBank[28][27] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[28][25]  ( .G(n17733), .D(n13250), .Q(\pipeline/RegFile_DEC_WB/RegBank[28][25] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[28][23]  ( .G(n17733), .D(n13244), .Q(\pipeline/RegFile_DEC_WB/RegBank[28][23] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[28][21]  ( .G(n13091), .D(n13238), .Q(\pipeline/RegFile_DEC_WB/RegBank[28][21] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[28][19]  ( .G(n17733), .D(n13232), .Q(\pipeline/RegFile_DEC_WB/RegBank[28][19] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[28][17]  ( .G(n13091), .D(n13226), .Q(\pipeline/RegFile_DEC_WB/RegBank[28][17] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[28][15]  ( .G(n17733), .D(n13220), .Q(\pipeline/RegFile_DEC_WB/RegBank[28][15] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[28][13]  ( .G(n13091), .D(n13214), .Q(\pipeline/RegFile_DEC_WB/RegBank[28][13] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[28][0]  ( .G(n17733), .D(n13175), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[28][0] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[28][8]  ( .G(n17733), .D(n13199), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[28][8] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[28][14]  ( .G(n13091), .D(n13217), .Q(\pipeline/RegFile_DEC_WB/RegBank[28][14] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[28][16]  ( .G(n17733), .D(n13223), .Q(\pipeline/RegFile_DEC_WB/RegBank[28][16] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[28][18]  ( .G(n17733), .D(n13229), .Q(\pipeline/RegFile_DEC_WB/RegBank[28][18] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[28][20]  ( .G(n13091), .D(n13235), .Q(\pipeline/RegFile_DEC_WB/RegBank[28][20] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[28][22]  ( .G(n13091), .D(n13241), .Q(\pipeline/RegFile_DEC_WB/RegBank[28][22] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[28][24]  ( .G(n13091), .D(n13247), .Q(\pipeline/RegFile_DEC_WB/RegBank[28][24] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[28][26]  ( .G(n13091), .D(n13253), .Q(\pipeline/RegFile_DEC_WB/RegBank[28][26] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[28][28]  ( .G(n13091), .D(n13259), .Q(\pipeline/RegFile_DEC_WB/RegBank[28][28] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[28][30]  ( .G(n17733), .D(n13265), .Q(\pipeline/RegFile_DEC_WB/RegBank[28][30] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[29][31]  ( .G(n13088), .D(n13268), .Q(\pipeline/RegFile_DEC_WB/RegBank[29][31] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[29][29]  ( .G(n17734), .D(n13262), .Q(\pipeline/RegFile_DEC_WB/RegBank[29][29] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[29][27]  ( .G(n13088), .D(n13256), .Q(\pipeline/RegFile_DEC_WB/RegBank[29][27] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[29][25]  ( .G(n17734), .D(n13250), .Q(\pipeline/RegFile_DEC_WB/RegBank[29][25] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[29][23]  ( .G(n17734), .D(n13244), .Q(\pipeline/RegFile_DEC_WB/RegBank[29][23] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[29][21]  ( .G(n13088), .D(n13238), .Q(\pipeline/RegFile_DEC_WB/RegBank[29][21] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[29][19]  ( .G(n17734), .D(n13232), .Q(\pipeline/RegFile_DEC_WB/RegBank[29][19] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[29][17]  ( .G(n13088), .D(n13226), .Q(\pipeline/RegFile_DEC_WB/RegBank[29][17] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[29][15]  ( .G(n17734), .D(n13220), .Q(\pipeline/RegFile_DEC_WB/RegBank[29][15] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[29][13]  ( .G(n13088), .D(n13214), .Q(\pipeline/RegFile_DEC_WB/RegBank[29][13] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[29][0]  ( .G(n17734), .D(n13175), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[29][0] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[29][8]  ( .G(n17734), .D(n13199), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[29][8] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[29][14]  ( .G(n13088), .D(n13217), .Q(\pipeline/RegFile_DEC_WB/RegBank[29][14] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[29][16]  ( .G(n17734), .D(n13223), .Q(\pipeline/RegFile_DEC_WB/RegBank[29][16] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[29][18]  ( .G(n17734), .D(n13229), .Q(\pipeline/RegFile_DEC_WB/RegBank[29][18] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[29][20]  ( .G(n13088), .D(n13235), .Q(\pipeline/RegFile_DEC_WB/RegBank[29][20] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[29][22]  ( .G(n13088), .D(n13241), .Q(\pipeline/RegFile_DEC_WB/RegBank[29][22] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[29][24]  ( .G(n13088), .D(n13247), .Q(\pipeline/RegFile_DEC_WB/RegBank[29][24] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[29][26]  ( .G(n13088), .D(n13253), .Q(\pipeline/RegFile_DEC_WB/RegBank[29][26] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[29][28]  ( .G(n13088), .D(n13259), .Q(\pipeline/RegFile_DEC_WB/RegBank[29][28] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[29][30]  ( .G(n17734), .D(n13265), .Q(\pipeline/RegFile_DEC_WB/RegBank[29][30] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[30][31]  ( .G(n13085), .D(n13268), .Q(\pipeline/RegFile_DEC_WB/RegBank[30][31] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[30][29]  ( .G(n17735), .D(n13262), .Q(\pipeline/RegFile_DEC_WB/RegBank[30][29] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[30][27]  ( .G(n13085), .D(n13256), .Q(\pipeline/RegFile_DEC_WB/RegBank[30][27] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[30][25]  ( .G(n17735), .D(n13250), .Q(\pipeline/RegFile_DEC_WB/RegBank[30][25] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[30][23]  ( .G(n17735), .D(n13244), .Q(\pipeline/RegFile_DEC_WB/RegBank[30][23] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[30][21]  ( .G(n13085), .D(n13238), .Q(\pipeline/RegFile_DEC_WB/RegBank[30][21] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[30][19]  ( .G(n17735), .D(n13232), .Q(\pipeline/RegFile_DEC_WB/RegBank[30][19] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[30][17]  ( .G(n13085), .D(n13226), .Q(\pipeline/RegFile_DEC_WB/RegBank[30][17] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[30][15]  ( .G(n17735), .D(n13220), .Q(\pipeline/RegFile_DEC_WB/RegBank[30][15] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[30][13]  ( .G(n13085), .D(n13214), .Q(\pipeline/RegFile_DEC_WB/RegBank[30][13] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[30][0]  ( .G(n17735), .D(n13175), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[30][0] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[30][8]  ( .G(n17735), .D(n13199), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[30][8] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[30][14]  ( .G(n13085), .D(n13217), .Q(\pipeline/RegFile_DEC_WB/RegBank[30][14] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[30][16]  ( .G(n17735), .D(n13223), .Q(\pipeline/RegFile_DEC_WB/RegBank[30][16] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[30][18]  ( .G(n17735), .D(n13229), .Q(\pipeline/RegFile_DEC_WB/RegBank[30][18] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[30][20]  ( .G(n13085), .D(n13235), .Q(\pipeline/RegFile_DEC_WB/RegBank[30][20] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[30][22]  ( .G(n13085), .D(n13241), .Q(\pipeline/RegFile_DEC_WB/RegBank[30][22] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[30][24]  ( .G(n13085), .D(n13247), .Q(\pipeline/RegFile_DEC_WB/RegBank[30][24] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[30][26]  ( .G(n13085), .D(n13253), .Q(\pipeline/RegFile_DEC_WB/RegBank[30][26] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[30][28]  ( .G(n13085), .D(n13259), .Q(\pipeline/RegFile_DEC_WB/RegBank[30][28] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[30][30]  ( .G(n17735), .D(n13265), .Q(\pipeline/RegFile_DEC_WB/RegBank[30][30] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[31][31]  ( .G(n13082), .D(n13268), .Q(\pipeline/RegFile_DEC_WB/RegBank[31][31] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg2_out_IDEX_reg[31]  ( .D(
        \pipeline/IDEX_Stage/N165 ), .CK(Clk), .Q(n13886), .QN(n17526) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[31][29]  ( .G(n17736), .D(n13262), .Q(\pipeline/RegFile_DEC_WB/RegBank[31][29] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg2_out_IDEX_reg[29]  ( .D(
        \pipeline/IDEX_Stage/N163 ), .CK(Clk), .Q(n13885), .QN(n17524) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[31][27]  ( .G(n13082), .D(n13256), .Q(\pipeline/RegFile_DEC_WB/RegBank[31][27] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg2_out_IDEX_reg[27]  ( .D(
        \pipeline/IDEX_Stage/N161 ), .CK(Clk), .Q(n13884), .QN(n17522) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[31][25]  ( .G(n17736), .D(n13250), .Q(\pipeline/RegFile_DEC_WB/RegBank[31][25] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg2_out_IDEX_reg[25]  ( .D(
        \pipeline/IDEX_Stage/N159 ), .CK(Clk), .Q(n13883), .QN(n17520) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[31][23]  ( .G(n17736), .D(n13244), .Q(\pipeline/RegFile_DEC_WB/RegBank[31][23] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg2_out_IDEX_reg[23]  ( .D(
        \pipeline/IDEX_Stage/N157 ), .CK(Clk), .Q(n13882), .QN(n17518) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[31][21]  ( .G(n13082), .D(n13238), .Q(\pipeline/RegFile_DEC_WB/RegBank[31][21] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg2_out_IDEX_reg[21]  ( .D(
        \pipeline/IDEX_Stage/N155 ), .CK(Clk), .Q(n13881), .QN(n17516) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[31][19]  ( .G(n17736), .D(n13232), .Q(\pipeline/RegFile_DEC_WB/RegBank[31][19] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg2_out_IDEX_reg[19]  ( .D(
        \pipeline/IDEX_Stage/N153 ), .CK(Clk), .Q(n13880), .QN(n17514) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[31][17]  ( .G(n13082), .D(n13226), .Q(\pipeline/RegFile_DEC_WB/RegBank[31][17] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg2_out_IDEX_reg[17]  ( .D(
        \pipeline/IDEX_Stage/N151 ), .CK(Clk), .Q(n13879), .QN(n17512) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[31][15]  ( .G(n17736), .D(n13220), .Q(\pipeline/RegFile_DEC_WB/RegBank[31][15] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg2_out_IDEX_reg[15]  ( .D(
        \pipeline/IDEX_Stage/N149 ), .CK(Clk), .Q(n13878), .QN(n17510) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[31][13]  ( .G(n13082), .D(n13214), .Q(\pipeline/RegFile_DEC_WB/RegBank[31][13] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg2_out_IDEX_reg[13]  ( .D(
        \pipeline/IDEX_Stage/N147 ), .CK(Clk), .Q(n13877), .QN(n17508) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[31][0]  ( .G(n17736), .D(n13175), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[31][0] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg2_out_IDEX_reg[0]  ( .D(
        \pipeline/IDEX_Stage/N134 ), .CK(Clk), .Q(n13876), .QN(n17495) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[31][8]  ( .G(n17736), .D(n13199), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[31][8] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg2_out_IDEX_reg[8]  ( .D(
        \pipeline/IDEX_Stage/N142 ), .CK(Clk), .Q(n13875), .QN(n17503) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[31][14]  ( .G(n13082), .D(n13217), .Q(\pipeline/RegFile_DEC_WB/RegBank[31][14] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg2_out_IDEX_reg[14]  ( .D(
        \pipeline/IDEX_Stage/N148 ), .CK(Clk), .Q(n13874), .QN(n17509) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[31][16]  ( .G(n17736), .D(n13223), .Q(\pipeline/RegFile_DEC_WB/RegBank[31][16] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg2_out_IDEX_reg[16]  ( .D(
        \pipeline/IDEX_Stage/N150 ), .CK(Clk), .Q(n13873), .QN(n17511) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[31][18]  ( .G(n17736), .D(n13229), .Q(\pipeline/RegFile_DEC_WB/RegBank[31][18] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg2_out_IDEX_reg[18]  ( .D(
        \pipeline/IDEX_Stage/N152 ), .CK(Clk), .Q(n13872), .QN(n17513) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[31][20]  ( .G(n13082), .D(n13235), .Q(\pipeline/RegFile_DEC_WB/RegBank[31][20] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg2_out_IDEX_reg[20]  ( .D(
        \pipeline/IDEX_Stage/N154 ), .CK(Clk), .Q(n13871), .QN(n17515) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[31][22]  ( .G(n13082), .D(n13241), .Q(\pipeline/RegFile_DEC_WB/RegBank[31][22] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg2_out_IDEX_reg[22]  ( .D(
        \pipeline/IDEX_Stage/N156 ), .CK(Clk), .Q(n13870), .QN(n17517) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[31][24]  ( .G(n13082), .D(n13247), .Q(\pipeline/RegFile_DEC_WB/RegBank[31][24] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg2_out_IDEX_reg[24]  ( .D(
        \pipeline/IDEX_Stage/N158 ), .CK(Clk), .Q(n13869), .QN(n17519) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[31][26]  ( .G(n13082), .D(n13253), .Q(\pipeline/RegFile_DEC_WB/RegBank[31][26] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg2_out_IDEX_reg[26]  ( .D(
        \pipeline/IDEX_Stage/N160 ), .CK(Clk), .Q(n13868), .QN(n17521) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[31][28]  ( .G(n13082), .D(n13259), .Q(\pipeline/RegFile_DEC_WB/RegBank[31][28] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg2_out_IDEX_reg[28]  ( .D(
        \pipeline/IDEX_Stage/N162 ), .CK(Clk), .Q(n13867), .QN(n17523) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[31][30]  ( .G(n17736), .D(n13265), .Q(\pipeline/RegFile_DEC_WB/RegBank[31][30] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg2_out_IDEX_reg[30]  ( .D(
        \pipeline/IDEX_Stage/N164 ), .CK(Clk), .Q(n13866), .QN(n17525) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_reg[28]  ( .D(n3912), .CK(Clk), .RN(
        n17705), .Q(n13865), .QN(n7675) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_reg[27]  ( .D(n3910), .CK(Clk), .RN(
        n17703), .Q(n13864), .QN(n7674) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_reg[26]  ( .D(n3908), .CK(Clk), .RN(
        n17702), .Q(n13863), .QN(n7673) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_reg[25]  ( .D(n3906), .CK(Clk), .RN(
        n17705), .Q(n13862), .QN(n7672) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_reg[24]  ( .D(n3904), .CK(Clk), .RN(
        n17705), .Q(n13861), .QN(n7671) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_reg[23]  ( .D(n3902), .CK(Clk), .RN(
        n17705), .Q(n13860), .QN(n7670) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_reg[22]  ( .D(n3900), .CK(Clk), .RN(
        n17703), .Q(n13859), .QN(n7669) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_reg[21]  ( .D(n3898), .CK(Clk), .RN(
        n17705), .Q(n13858), .QN(n7668) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_reg[20]  ( .D(n3896), .CK(Clk), .RN(
        n17705), .Q(n13857), .QN(n7667) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_reg[19]  ( .D(n3894), .CK(Clk), .RN(
        n17704), .Q(n13856), .QN(n7666) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_reg[18]  ( .D(n3892), .CK(Clk), .RN(
        n17705), .Q(n13855), .QN(n7665) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_reg[17]  ( .D(n3890), .CK(Clk), .RN(
        n17705), .Q(n13854), .QN(n7664) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_reg[15]  ( .D(n3888), .CK(Clk), .RN(
        n17705), .Q(n13853), .QN(n7663) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_reg[14]  ( .D(n3886), .CK(Clk), .RN(
        n17705), .Q(n13852), .QN(n7662) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_reg[13]  ( .D(n3884), .CK(Clk), .RN(
        n17701), .Q(n13851), .QN(n7661) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_reg[8]  ( .D(n3882), .CK(Clk), .RN(
        n17705), .Q(n13850), .QN(n7660) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_reg[0]  ( .D(n3880), .CK(Clk), .RN(
        n17704), .Q(n13849), .QN(n7659) );
  DLH_X1 \DataMem/Mem_reg[0][1]  ( .G(n13058), .D(\DataMem/N1651 ), .Q(
        \DataMem/Mem[0][1] ) );
  DLL_X1 \DataMem/Dataout_reg[1]  ( .D(\DataMem/N2164 ), .GN(n17098), .Q(
        \DataMem/N2346 ) );
  DFF_X1 \pipeline/MEMWB_Stage/Data_to_RF_reg[1]  ( .D(
        \pipeline/MEMWB_Stage/N12 ), .CK(Clk), .Q(
        \pipeline/data_to_RF_from_WB[1] ), .QN(n17321) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[2][1]  ( .G(n17707), .D(n13178), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[2][1] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[4][1]  ( .G(n17709), .D(n13178), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[4][1] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[6][1]  ( .G(n17711), .D(n13178), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[6][1] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[8][1]  ( .G(n17713), .D(n13178), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[8][1] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[10][1]  ( .G(n17715), .D(n13178), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[10][1] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[12][1]  ( .G(n17717), .D(n13178), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[12][1] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[14][1]  ( .G(n17719), .D(n13178), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[14][1] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[16][1]  ( .G(n17721), .D(n13178), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[16][1] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[18][1]  ( .G(n17723), .D(n13178), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[18][1] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[20][1]  ( .G(n17725), .D(n13178), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[20][1] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[22][1]  ( .G(n17727), .D(n13178), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[22][1] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[24][1]  ( .G(n17729), .D(n13178), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[24][1] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[26][1]  ( .G(n17731), .D(n13178), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[26][1] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[28][1]  ( .G(n17733), .D(n13178), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[28][1] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[30][1]  ( .G(n17735), .D(n13178), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[30][1] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[31][1]  ( .G(n17736), .D(n13178), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[31][1] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[29][1]  ( .G(n17734), .D(n13178), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[29][1] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[27][1]  ( .G(n17732), .D(n13178), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[27][1] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[25][1]  ( .G(n17730), .D(n13178), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[25][1] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[23][1]  ( .G(n17728), .D(n13178), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[23][1] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[21][1]  ( .G(n17726), .D(n13178), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[21][1] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[19][1]  ( .G(n17724), .D(n13178), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[19][1] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[17][1]  ( .G(n17722), .D(n13178), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[17][1] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[15][1]  ( .G(n17720), .D(n13178), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[15][1] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[13][1]  ( .G(n17718), .D(n13178), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[13][1] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[11][1]  ( .G(n17716), .D(n13178), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[11][1] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[9][1]  ( .G(n17714), .D(n13178), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[9][1] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[7][1]  ( .G(n17712), .D(n13178), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[7][1] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[5][1]  ( .G(n17710), .D(n13178), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[5][1] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[3][1]  ( .G(n17708), .D(n13178), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[3][1] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[1][1]  ( .G(n17706), .D(n13178), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[1][1] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg2_out_IDEX_reg[1]  ( .D(
        \pipeline/IDEX_Stage/N135 ), .CK(Clk), .Q(n13848), .QN(n17496) );
  DFF_X1 \pipeline/IDEX_Stage/Reg1_out_IDEX_reg[1]  ( .D(
        \pipeline/IDEX_Stage/N103 ), .CK(Clk), .Q(n13847) );
  DFF_X1 \pipeline/MEMWB_Stage/Data_to_RF_reg[3]  ( .D(
        \pipeline/MEMWB_Stage/N14 ), .CK(Clk), .Q(
        \pipeline/data_to_RF_from_WB[3] ), .QN(n17306) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[2][3]  ( .G(n17707), .D(n13184), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[2][3] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[4][3]  ( .G(n17709), .D(n13184), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[4][3] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[6][3]  ( .G(n17711), .D(n13184), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[6][3] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[8][3]  ( .G(n17713), .D(n13184), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[8][3] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[10][3]  ( .G(n17715), .D(n13184), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[10][3] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[12][3]  ( .G(n17717), .D(n13184), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[12][3] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[14][3]  ( .G(n17719), .D(n13184), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[14][3] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[16][3]  ( .G(n17721), .D(n13184), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[16][3] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[18][3]  ( .G(n17723), .D(n13184), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[18][3] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[20][3]  ( .G(n17725), .D(n13184), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[20][3] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[22][3]  ( .G(n17727), .D(n13184), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[22][3] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[24][3]  ( .G(n17729), .D(n13184), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[24][3] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[26][3]  ( .G(n17731), .D(n13184), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[26][3] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[28][3]  ( .G(n17733), .D(n13184), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[28][3] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[30][3]  ( .G(n17735), .D(n13184), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[30][3] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[31][3]  ( .G(n17736), .D(n13184), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[31][3] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[29][3]  ( .G(n17734), .D(n13184), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[29][3] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[27][3]  ( .G(n17732), .D(n13184), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[27][3] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[25][3]  ( .G(n17730), .D(n13184), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[25][3] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[23][3]  ( .G(n17728), .D(n13184), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[23][3] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[21][3]  ( .G(n17726), .D(n13184), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[21][3] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[19][3]  ( .G(n17724), .D(n13184), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[19][3] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[17][3]  ( .G(n17722), .D(n13184), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[17][3] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[15][3]  ( .G(n17720), .D(n13184), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[15][3] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[13][3]  ( .G(n17718), .D(n13184), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[13][3] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[11][3]  ( .G(n17716), .D(n13184), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[11][3] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[9][3]  ( .G(n17714), .D(n13184), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[9][3] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[7][3]  ( .G(n17712), .D(n13184), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[7][3] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[5][3]  ( .G(n17710), .D(n13184), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[5][3] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[3][3]  ( .G(n17708), .D(n13184), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[3][3] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[1][3]  ( .G(n17706), .D(n13184), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[1][3] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg2_out_IDEX_reg[3]  ( .D(
        \pipeline/IDEX_Stage/N137 ), .CK(Clk), .Q(n13846), .QN(n17498) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_reg[3]  ( .D(n3878), .CK(Clk), .RN(
        n17704), .Q(n13845), .QN(n7658) );
  DFF_X1 \pipeline/IDEX_Stage/Reg1_out_IDEX_reg[3]  ( .D(
        \pipeline/IDEX_Stage/N105 ), .CK(Clk), .Q(n13844) );
  DLH_X1 \DataMem/Mem_reg[0][6]  ( .G(n13058), .D(\DataMem/N1661 ), .Q(
        \DataMem/Mem[0][6] ) );
  DLL_X1 \DataMem/Dataout_reg[6]  ( .D(\DataMem/N2179 ), .GN(n17098), .Q(
        \DataMem/N2331 ) );
  DFF_X1 \pipeline/MEMWB_Stage/Data_to_RF_reg[6]  ( .D(
        \pipeline/MEMWB_Stage/N17 ), .CK(Clk), .Q(
        \pipeline/data_to_RF_from_WB[6] ), .QN(n17318) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[2][6]  ( .G(n17707), .D(n13193), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[2][6] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[4][6]  ( .G(n17709), .D(n13193), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[4][6] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[6][6]  ( .G(n17711), .D(n13193), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[6][6] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[8][6]  ( .G(n17713), .D(n13193), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[8][6] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[10][6]  ( .G(n17715), .D(n13193), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[10][6] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[12][6]  ( .G(n17717), .D(n13193), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[12][6] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[14][6]  ( .G(n17719), .D(n13193), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[14][6] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[16][6]  ( .G(n17721), .D(n13193), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[16][6] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[18][6]  ( .G(n17723), .D(n13193), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[18][6] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[20][6]  ( .G(n17725), .D(n13193), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[20][6] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[22][6]  ( .G(n17727), .D(n13193), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[22][6] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[24][6]  ( .G(n17729), .D(n13193), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[24][6] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[26][6]  ( .G(n17731), .D(n13193), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[26][6] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[28][6]  ( .G(n17733), .D(n13193), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[28][6] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[30][6]  ( .G(n17735), .D(n13193), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[30][6] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[31][6]  ( .G(n17736), .D(n13193), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[31][6] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[29][6]  ( .G(n17734), .D(n13193), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[29][6] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[27][6]  ( .G(n17732), .D(n13193), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[27][6] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[25][6]  ( .G(n17730), .D(n13193), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[25][6] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[23][6]  ( .G(n17728), .D(n13193), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[23][6] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[21][6]  ( .G(n17726), .D(n13193), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[21][6] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[19][6]  ( .G(n17724), .D(n13193), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[19][6] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[17][6]  ( .G(n17722), .D(n13193), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[17][6] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[15][6]  ( .G(n17720), .D(n13193), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[15][6] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[13][6]  ( .G(n17718), .D(n13193), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[13][6] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[11][6]  ( .G(n17716), .D(n13193), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[11][6] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[9][6]  ( .G(n17714), .D(n13193), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[9][6] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[7][6]  ( .G(n17712), .D(n13193), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[7][6] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[5][6]  ( .G(n17710), .D(n13193), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[5][6] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[3][6]  ( .G(n17708), .D(n13193), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[3][6] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[1][6]  ( .G(n17706), .D(n13193), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[1][6] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg2_out_IDEX_reg[6]  ( .D(
        \pipeline/IDEX_Stage/N140 ), .CK(Clk), .Q(n13843), .QN(n17501) );
  DFF_X1 \pipeline/IDEX_Stage/Reg1_out_IDEX_reg[6]  ( .D(
        \pipeline/IDEX_Stage/N108 ), .CK(Clk), .Q(n13842) );
  DFF_X1 \pipeline/EXMEM_stage/ALUres_MEMaddr_out_EXMEM_reg[7]  ( .D(
        \pipeline/EXMEM_stage/N14 ), .CK(Clk), .Q(
        \pipeline/Alu_Out_Addr_to_mem[7] ) );
  DFF_X1 \pipeline/MEMWB_Stage/Data_to_RF_reg[7]  ( .D(
        \pipeline/MEMWB_Stage/N18 ), .CK(Clk), .Q(
        \pipeline/data_to_RF_from_WB[7] ), .QN(n17343) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[2][7]  ( .G(n17707), .D(n13196), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[2][7] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[4][7]  ( .G(n17709), .D(n13196), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[4][7] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[6][7]  ( .G(n17711), .D(n13196), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[6][7] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[8][7]  ( .G(n17713), .D(n13196), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[8][7] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[10][7]  ( .G(n17715), .D(n13196), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[10][7] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[12][7]  ( .G(n17717), .D(n13196), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[12][7] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[14][7]  ( .G(n17719), .D(n13196), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[14][7] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[16][7]  ( .G(n17721), .D(n13196), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[16][7] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[18][7]  ( .G(n17723), .D(n13196), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[18][7] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[20][7]  ( .G(n17725), .D(n13196), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[20][7] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[22][7]  ( .G(n17727), .D(n13196), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[22][7] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[24][7]  ( .G(n17729), .D(n13196), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[24][7] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[26][7]  ( .G(n17731), .D(n13196), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[26][7] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[28][7]  ( .G(n17733), .D(n13196), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[28][7] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[30][7]  ( .G(n17735), .D(n13196), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[30][7] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[31][7]  ( .G(n17736), .D(n13196), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[31][7] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[29][7]  ( .G(n17734), .D(n13196), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[29][7] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[27][7]  ( .G(n17732), .D(n13196), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[27][7] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[25][7]  ( .G(n17730), .D(n13196), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[25][7] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[23][7]  ( .G(n17728), .D(n13196), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[23][7] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[21][7]  ( .G(n17726), .D(n13196), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[21][7] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[19][7]  ( .G(n17724), .D(n13196), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[19][7] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[17][7]  ( .G(n17722), .D(n13196), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[17][7] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[15][7]  ( .G(n17720), .D(n13196), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[15][7] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[13][7]  ( .G(n17718), .D(n13196), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[13][7] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[11][7]  ( .G(n17716), .D(n13196), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[11][7] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[9][7]  ( .G(n17714), .D(n13196), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[9][7] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[7][7]  ( .G(n17712), .D(n13196), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[7][7] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[5][7]  ( .G(n17710), .D(n13196), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[5][7] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[3][7]  ( .G(n17708), .D(n13196), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[3][7] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[1][7]  ( .G(n17706), .D(n13196), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[1][7] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg2_out_IDEX_reg[7]  ( .D(
        \pipeline/IDEX_Stage/N141 ), .CK(Clk), .Q(n13841), .QN(n17502) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_reg[7]  ( .D(n3876), .CK(Clk), .RN(
        n17705), .Q(n13840), .QN(n7657) );
  DFF_X1 \pipeline/IDEX_Stage/Reg1_out_IDEX_reg[7]  ( .D(
        \pipeline/IDEX_Stage/N109 ), .CK(Clk), .Q(n13839) );
  DLH_X1 \DataMem/Mem_reg[7][1]  ( .G(n13079), .D(\DataMem/N2099 ), .Q(
        \DataMem/Mem[7][1] ) );
  DLH_X1 \DataMem/Mem_reg[6][1]  ( .G(n13076), .D(\DataMem/N2035 ), .Q(
        \DataMem/Mem[6][1] ) );
  DLH_X1 \DataMem/Mem_reg[5][1]  ( .G(n13073), .D(\DataMem/N1971 ), .Q(
        \DataMem/Mem[5][1] ) );
  DLH_X1 \DataMem/Mem_reg[4][1]  ( .G(n13070), .D(\DataMem/N1907 ), .Q(
        \DataMem/Mem[4][1] ) );
  DLH_X1 \DataMem/Mem_reg[3][1]  ( .G(n13067), .D(\DataMem/N1843 ), .Q(
        \DataMem/Mem[3][1] ) );
  DLH_X1 \DataMem/Mem_reg[2][1]  ( .G(n13064), .D(\DataMem/N1779 ), .Q(
        \DataMem/Mem[2][1] ) );
  DLH_X1 \DataMem/Mem_reg[1][1]  ( .G(n13061), .D(\DataMem/N1715 ), .Q(
        \DataMem/Mem[1][1] ) );
  DFF_X1 \pipeline/MEMWB_Stage/Data_to_RF_reg[4]  ( .D(
        \pipeline/MEMWB_Stage/N15 ), .CK(Clk), .Q(
        \pipeline/data_to_RF_from_WB[4] ), .QN(n17320) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[2][4]  ( .G(n17707), .D(n13187), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[2][4] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[4][4]  ( .G(n17709), .D(n13187), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[4][4] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[6][4]  ( .G(n17711), .D(n13187), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[6][4] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[8][4]  ( .G(n17713), .D(n13187), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[8][4] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[10][4]  ( .G(n17715), .D(n13187), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[10][4] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[12][4]  ( .G(n17717), .D(n13187), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[12][4] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[14][4]  ( .G(n17719), .D(n13187), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[14][4] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[16][4]  ( .G(n17721), .D(n13187), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[16][4] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[18][4]  ( .G(n17723), .D(n13187), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[18][4] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[20][4]  ( .G(n17725), .D(n13187), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[20][4] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[22][4]  ( .G(n17727), .D(n13187), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[22][4] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[24][4]  ( .G(n17729), .D(n13187), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[24][4] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[26][4]  ( .G(n17731), .D(n13187), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[26][4] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[28][4]  ( .G(n17733), .D(n13187), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[28][4] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[30][4]  ( .G(n17735), .D(n13187), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[30][4] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[31][4]  ( .G(n17736), .D(n13187), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[31][4] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[29][4]  ( .G(n17734), .D(n13187), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[29][4] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[27][4]  ( .G(n17732), .D(n13187), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[27][4] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[25][4]  ( .G(n17730), .D(n13187), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[25][4] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[23][4]  ( .G(n17728), .D(n13187), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[23][4] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[21][4]  ( .G(n17726), .D(n13187), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[21][4] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[19][4]  ( .G(n17724), .D(n13187), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[19][4] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[17][4]  ( .G(n17722), .D(n13187), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[17][4] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[15][4]  ( .G(n17720), .D(n13187), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[15][4] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[13][4]  ( .G(n17718), .D(n13187), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[13][4] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[11][4]  ( .G(n17716), .D(n13187), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[11][4] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[9][4]  ( .G(n17714), .D(n13187), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[9][4] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[7][4]  ( .G(n17712), .D(n13187), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[7][4] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[5][4]  ( .G(n17710), .D(n13187), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[5][4] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[3][4]  ( .G(n17708), .D(n13187), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[3][4] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[1][4]  ( .G(n17706), .D(n13187), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[1][4] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg2_out_IDEX_reg[4]  ( .D(
        \pipeline/IDEX_Stage/N138 ), .CK(Clk), .Q(n13838), .QN(n17499) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_reg[4]  ( .D(n3874), .CK(Clk), .RN(
        n17704), .Q(n13837), .QN(n7656) );
  DFF_X1 \pipeline/IDEX_Stage/Reg1_out_IDEX_reg[4]  ( .D(
        \pipeline/IDEX_Stage/N106 ), .CK(Clk), .Q(n13836) );
  DFF_X1 \pipeline/EXMEM_stage/DataToMem_out_EXMEM_reg[4]  ( .D(
        \pipeline/EXMEM_stage/N43 ), .CK(Clk), .Q(n13835) );
  DLH_X1 \DataMem/Mem_reg[7][4]  ( .G(n13079), .D(\DataMem/N2105 ), .Q(
        \DataMem/Mem[7][4] ) );
  DLH_X1 \DataMem/Mem_reg[6][4]  ( .G(n13076), .D(\DataMem/N2041 ), .Q(
        \DataMem/Mem[6][4] ) );
  DLH_X1 \DataMem/Mem_reg[5][4]  ( .G(n13073), .D(\DataMem/N1977 ), .Q(
        \DataMem/Mem[5][4] ) );
  DLH_X1 \DataMem/Mem_reg[4][4]  ( .G(n13070), .D(\DataMem/N1913 ), .Q(
        \DataMem/Mem[4][4] ) );
  DLH_X1 \DataMem/Mem_reg[3][4]  ( .G(n13067), .D(\DataMem/N1849 ), .Q(
        \DataMem/Mem[3][4] ) );
  DLH_X1 \DataMem/Mem_reg[2][4]  ( .G(n13064), .D(\DataMem/N1785 ), .Q(
        \DataMem/Mem[2][4] ) );
  DLH_X1 \DataMem/Mem_reg[1][4]  ( .G(n13061), .D(\DataMem/N1721 ), .Q(
        \DataMem/Mem[1][4] ) );
  DLH_X1 \DataMem/Mem_reg[0][4]  ( .G(n13058), .D(\DataMem/N1657 ), .Q(
        \DataMem/Mem[0][4] ) );
  DLL_X1 \DataMem/Dataout_reg[4]  ( .D(\DataMem/N2173 ), .GN(n17098), .Q(
        \DataMem/N2337 ) );
  DFF_X1 \pipeline/MEMWB_Stage/Data_to_RF_reg[5]  ( .D(
        \pipeline/MEMWB_Stage/N16 ), .CK(Clk), .Q(
        \pipeline/data_to_RF_from_WB[5] ), .QN(n17308) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[2][5]  ( .G(n13169), .D(n13190), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[2][5] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[4][5]  ( .G(n13163), .D(n13190), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[4][5] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[6][5]  ( .G(n13157), .D(n13190), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[6][5] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[8][5]  ( .G(n13151), .D(n13190), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[8][5] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[10][5]  ( .G(n13145), .D(n13190), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[10][5] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[12][5]  ( .G(n13139), .D(n13190), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[12][5] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[14][5]  ( .G(n13133), .D(n13190), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[14][5] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[16][5]  ( .G(n13127), .D(n13190), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[16][5] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[18][5]  ( .G(n13121), .D(n13190), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[18][5] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[20][5]  ( .G(n13115), .D(n13190), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[20][5] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[22][5]  ( .G(n13109), .D(n13190), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[22][5] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[24][5]  ( .G(n13103), .D(n13190), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[24][5] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[26][5]  ( .G(n13097), .D(n13190), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[26][5] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[28][5]  ( .G(n13091), .D(n13190), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[28][5] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[30][5]  ( .G(n13085), .D(n13190), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[30][5] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[31][5]  ( .G(n13082), .D(n13190), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[31][5] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[29][5]  ( .G(n13088), .D(n13190), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[29][5] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[27][5]  ( .G(n13094), .D(n13190), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[27][5] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[25][5]  ( .G(n13100), .D(n13190), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[25][5] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[23][5]  ( .G(n13106), .D(n13190), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[23][5] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[21][5]  ( .G(n13112), .D(n13190), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[21][5] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[19][5]  ( .G(n13118), .D(n13190), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[19][5] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[17][5]  ( .G(n13124), .D(n13190), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[17][5] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[15][5]  ( .G(n13130), .D(n13190), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[15][5] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[13][5]  ( .G(n13136), .D(n13190), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[13][5] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[11][5]  ( .G(n13142), .D(n13190), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[11][5] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[9][5]  ( .G(n13148), .D(n13190), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[9][5] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[7][5]  ( .G(n13154), .D(n13190), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[7][5] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[5][5]  ( .G(n13160), .D(n13190), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[5][5] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[3][5]  ( .G(n13166), .D(n13190), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[3][5] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[1][5]  ( .G(n13172), .D(n13190), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[1][5] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg2_out_IDEX_reg[5]  ( .D(
        \pipeline/IDEX_Stage/N139 ), .CK(Clk), .Q(n13834), .QN(n17500) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_reg[5]  ( .D(n3872), .CK(Clk), .RN(
        n17705), .Q(n13833), .QN(n7655) );
  DFF_X1 \pipeline/IDEX_Stage/Reg1_out_IDEX_reg[5]  ( .D(
        \pipeline/IDEX_Stage/N107 ), .CK(Clk), .Q(n13832) );
  DFF_X1 \pipeline/EXMEM_stage/DataToMem_out_EXMEM_reg[5]  ( .D(
        \pipeline/EXMEM_stage/N44 ), .CK(Clk), .Q(n13831) );
  DLH_X1 \DataMem/Mem_reg[7][5]  ( .G(n13079), .D(\DataMem/N2107 ), .Q(
        \DataMem/Mem[7][5] ) );
  DLH_X1 \DataMem/Mem_reg[6][5]  ( .G(n13076), .D(\DataMem/N2043 ), .Q(
        \DataMem/Mem[6][5] ) );
  DLH_X1 \DataMem/Mem_reg[5][5]  ( .G(n13073), .D(\DataMem/N1979 ), .Q(
        \DataMem/Mem[5][5] ) );
  DLH_X1 \DataMem/Mem_reg[4][5]  ( .G(n13070), .D(\DataMem/N1915 ), .Q(
        \DataMem/Mem[4][5] ) );
  DLH_X1 \DataMem/Mem_reg[3][5]  ( .G(n13067), .D(\DataMem/N1851 ), .Q(
        \DataMem/Mem[3][5] ) );
  DLH_X1 \DataMem/Mem_reg[2][5]  ( .G(n13064), .D(\DataMem/N1787 ), .Q(
        \DataMem/Mem[2][5] ) );
  DLH_X1 \DataMem/Mem_reg[1][5]  ( .G(n13061), .D(\DataMem/N1723 ), .Q(
        \DataMem/Mem[1][5] ) );
  DLH_X1 \DataMem/Mem_reg[0][5]  ( .G(n13058), .D(\DataMem/N1659 ), .Q(
        \DataMem/Mem[0][5] ) );
  DLL_X1 \DataMem/Dataout_reg[5]  ( .D(\DataMem/N2176 ), .GN(n17098), .Q(
        \DataMem/N2334 ) );
  DFF_X1 \pipeline/EXMEM_stage/DataToMem_out_EXMEM_reg[7]  ( .D(
        \pipeline/EXMEM_stage/N46 ), .CK(Clk), .Q(n13830) );
  DLH_X1 \DataMem/Mem_reg[7][7]  ( .G(n13079), .D(\DataMem/N2111 ), .Q(
        \DataMem/Mem[7][7] ) );
  DLH_X1 \DataMem/Mem_reg[6][7]  ( .G(n13076), .D(\DataMem/N2047 ), .Q(
        \DataMem/Mem[6][7] ) );
  DLH_X1 \DataMem/Mem_reg[5][7]  ( .G(n13073), .D(\DataMem/N1983 ), .Q(
        \DataMem/Mem[5][7] ) );
  DLH_X1 \DataMem/Mem_reg[4][7]  ( .G(n13070), .D(\DataMem/N1919 ), .Q(
        \DataMem/Mem[4][7] ) );
  DLH_X1 \DataMem/Mem_reg[3][7]  ( .G(n13067), .D(\DataMem/N1855 ), .Q(
        \DataMem/Mem[3][7] ) );
  DLH_X1 \DataMem/Mem_reg[2][7]  ( .G(n13064), .D(\DataMem/N1791 ), .Q(
        \DataMem/Mem[2][7] ) );
  DLH_X1 \DataMem/Mem_reg[1][7]  ( .G(n13061), .D(\DataMem/N1727 ), .Q(
        \DataMem/Mem[1][7] ) );
  DLH_X1 \DataMem/Mem_reg[0][7]  ( .G(n13058), .D(\DataMem/N1663 ), .Q(
        \DataMem/Mem[0][7] ) );
  DLL_X1 \DataMem/Dataout_reg[7]  ( .D(\DataMem/N2182 ), .GN(n17098), .Q(
        \DataMem/N2328 ) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_reg[6]  ( .D(n3870), .CK(Clk), .RN(
        n17705), .Q(n13829), .QN(n7654) );
  DFF_X1 \pipeline/EXMEM_stage/DataToMem_out_EXMEM_reg[6]  ( .D(
        \pipeline/EXMEM_stage/N45 ), .CK(Clk), .Q(n13828) );
  DLH_X1 \DataMem/Mem_reg[7][6]  ( .G(n13079), .D(\DataMem/N2109 ), .Q(
        \DataMem/Mem[7][6] ) );
  DLH_X1 \DataMem/Mem_reg[6][6]  ( .G(n13076), .D(\DataMem/N2045 ), .Q(
        \DataMem/Mem[6][6] ) );
  DLH_X1 \DataMem/Mem_reg[5][6]  ( .G(n13073), .D(\DataMem/N1981 ), .Q(
        \DataMem/Mem[5][6] ) );
  DLH_X1 \DataMem/Mem_reg[4][6]  ( .G(n13070), .D(\DataMem/N1917 ), .Q(
        \DataMem/Mem[4][6] ) );
  DLH_X1 \DataMem/Mem_reg[3][6]  ( .G(n13067), .D(\DataMem/N1853 ), .Q(
        \DataMem/Mem[3][6] ) );
  DLH_X1 \DataMem/Mem_reg[2][6]  ( .G(n13064), .D(\DataMem/N1789 ), .Q(
        \DataMem/Mem[2][6] ) );
  DLH_X1 \DataMem/Mem_reg[1][6]  ( .G(n13061), .D(\DataMem/N1725 ), .Q(
        \DataMem/Mem[1][6] ) );
  DLH_X1 \DataMem/Mem_reg[0][10]  ( .G(n13058), .D(\DataMem/N1669 ), .Q(
        \DataMem/Mem[0][10] ) );
  DLL_X1 \DataMem/Dataout_reg[10]  ( .D(\DataMem/N2191 ), .GN(n13055), .Q(
        \DataMem/N2319 ) );
  DFF_X1 \pipeline/MEMWB_Stage/Data_to_RF_reg[10]  ( .D(
        \pipeline/MEMWB_Stage/N21 ), .CK(Clk), .Q(
        \pipeline/data_to_RF_from_WB[10] ), .QN(n17307) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[2][10]  ( .G(n13169), .D(n13205), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[2][10] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[4][10]  ( .G(n13163), .D(n13205), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[4][10] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[6][10]  ( .G(n13157), .D(n13205), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[6][10] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[8][10]  ( .G(n13151), .D(n13205), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[8][10] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[10][10]  ( .G(n13145), .D(n13205), .Q(\pipeline/RegFile_DEC_WB/RegBank[10][10] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[12][10]  ( .G(n13139), .D(n13205), .Q(\pipeline/RegFile_DEC_WB/RegBank[12][10] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[14][10]  ( .G(n13133), .D(n13205), .Q(\pipeline/RegFile_DEC_WB/RegBank[14][10] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[16][10]  ( .G(n13127), .D(n13205), .Q(\pipeline/RegFile_DEC_WB/RegBank[16][10] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[18][10]  ( .G(n13121), .D(n13205), .Q(\pipeline/RegFile_DEC_WB/RegBank[18][10] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[20][10]  ( .G(n13115), .D(n13205), .Q(\pipeline/RegFile_DEC_WB/RegBank[20][10] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[22][10]  ( .G(n13109), .D(n13205), .Q(\pipeline/RegFile_DEC_WB/RegBank[22][10] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[24][10]  ( .G(n13103), .D(n13205), .Q(\pipeline/RegFile_DEC_WB/RegBank[24][10] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[26][10]  ( .G(n13097), .D(n13205), .Q(\pipeline/RegFile_DEC_WB/RegBank[26][10] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[28][10]  ( .G(n13091), .D(n13205), .Q(\pipeline/RegFile_DEC_WB/RegBank[28][10] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[30][10]  ( .G(n13085), .D(n13205), .Q(\pipeline/RegFile_DEC_WB/RegBank[30][10] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[31][10]  ( .G(n13082), .D(n13205), .Q(\pipeline/RegFile_DEC_WB/RegBank[31][10] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[29][10]  ( .G(n13088), .D(n13205), .Q(\pipeline/RegFile_DEC_WB/RegBank[29][10] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[27][10]  ( .G(n13094), .D(n13205), .Q(\pipeline/RegFile_DEC_WB/RegBank[27][10] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[25][10]  ( .G(n13100), .D(n13205), .Q(\pipeline/RegFile_DEC_WB/RegBank[25][10] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[23][10]  ( .G(n13106), .D(n13205), .Q(\pipeline/RegFile_DEC_WB/RegBank[23][10] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[21][10]  ( .G(n13112), .D(n13205), .Q(\pipeline/RegFile_DEC_WB/RegBank[21][10] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[19][10]  ( .G(n13118), .D(n13205), .Q(\pipeline/RegFile_DEC_WB/RegBank[19][10] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[17][10]  ( .G(n13124), .D(n13205), .Q(\pipeline/RegFile_DEC_WB/RegBank[17][10] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[15][10]  ( .G(n13130), .D(n13205), .Q(\pipeline/RegFile_DEC_WB/RegBank[15][10] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[13][10]  ( .G(n13136), .D(n13205), .Q(\pipeline/RegFile_DEC_WB/RegBank[13][10] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[11][10]  ( .G(n13142), .D(n13205), .Q(\pipeline/RegFile_DEC_WB/RegBank[11][10] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[9][10]  ( .G(n13148), .D(n13205), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[9][10] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[7][10]  ( .G(n13154), .D(n13205), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[7][10] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[5][10]  ( .G(n13160), .D(n13205), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[5][10] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[3][10]  ( .G(n13166), .D(n13205), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[3][10] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[1][10]  ( .G(n13172), .D(n13205), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[1][10] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg2_out_IDEX_reg[10]  ( .D(
        \pipeline/IDEX_Stage/N144 ), .CK(Clk), .Q(n13827), .QN(n17505) );
  DFF_X1 \pipeline/IDEX_Stage/Reg1_out_IDEX_reg[10]  ( .D(
        \pipeline/IDEX_Stage/N112 ), .CK(Clk), .Q(n13826) );
  DFF_X1 \pipeline/MEMWB_Stage/Data_to_RF_reg[11]  ( .D(
        \pipeline/MEMWB_Stage/N22 ), .CK(Clk), .Q(
        \pipeline/data_to_RF_from_WB[11] ), .QN(n17319) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[2][11]  ( .G(n17707), .D(n13208), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[2][11] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[4][11]  ( .G(n17709), .D(n13208), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[4][11] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[6][11]  ( .G(n17711), .D(n13208), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[6][11] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[8][11]  ( .G(n17713), .D(n13208), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[8][11] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[10][11]  ( .G(n17715), .D(n13208), .Q(\pipeline/RegFile_DEC_WB/RegBank[10][11] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[12][11]  ( .G(n17717), .D(n13208), .Q(\pipeline/RegFile_DEC_WB/RegBank[12][11] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[14][11]  ( .G(n17719), .D(n13208), .Q(\pipeline/RegFile_DEC_WB/RegBank[14][11] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[16][11]  ( .G(n17721), .D(n13208), .Q(\pipeline/RegFile_DEC_WB/RegBank[16][11] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[18][11]  ( .G(n17723), .D(n13208), .Q(\pipeline/RegFile_DEC_WB/RegBank[18][11] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[20][11]  ( .G(n17725), .D(n13208), .Q(\pipeline/RegFile_DEC_WB/RegBank[20][11] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[22][11]  ( .G(n17727), .D(n13208), .Q(\pipeline/RegFile_DEC_WB/RegBank[22][11] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[24][11]  ( .G(n17729), .D(n13208), .Q(\pipeline/RegFile_DEC_WB/RegBank[24][11] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[26][11]  ( .G(n17731), .D(n13208), .Q(\pipeline/RegFile_DEC_WB/RegBank[26][11] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[28][11]  ( .G(n17733), .D(n13208), .Q(\pipeline/RegFile_DEC_WB/RegBank[28][11] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[30][11]  ( .G(n17735), .D(n13208), .Q(\pipeline/RegFile_DEC_WB/RegBank[30][11] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[31][11]  ( .G(n17736), .D(n13208), .Q(\pipeline/RegFile_DEC_WB/RegBank[31][11] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[29][11]  ( .G(n17734), .D(n13208), .Q(\pipeline/RegFile_DEC_WB/RegBank[29][11] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[27][11]  ( .G(n17732), .D(n13208), .Q(\pipeline/RegFile_DEC_WB/RegBank[27][11] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[25][11]  ( .G(n17730), .D(n13208), .Q(\pipeline/RegFile_DEC_WB/RegBank[25][11] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[23][11]  ( .G(n17728), .D(n13208), .Q(\pipeline/RegFile_DEC_WB/RegBank[23][11] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[21][11]  ( .G(n17726), .D(n13208), .Q(\pipeline/RegFile_DEC_WB/RegBank[21][11] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[19][11]  ( .G(n17724), .D(n13208), .Q(\pipeline/RegFile_DEC_WB/RegBank[19][11] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[17][11]  ( .G(n17722), .D(n13208), .Q(\pipeline/RegFile_DEC_WB/RegBank[17][11] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[15][11]  ( .G(n17720), .D(n13208), .Q(\pipeline/RegFile_DEC_WB/RegBank[15][11] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[13][11]  ( .G(n17718), .D(n13208), .Q(\pipeline/RegFile_DEC_WB/RegBank[13][11] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[11][11]  ( .G(n17716), .D(n13208), .Q(\pipeline/RegFile_DEC_WB/RegBank[11][11] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[9][11]  ( .G(n17714), .D(n13208), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[9][11] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[7][11]  ( .G(n17712), .D(n13208), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[7][11] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[5][11]  ( .G(n17710), .D(n13208), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[5][11] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[3][11]  ( .G(n17708), .D(n13208), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[3][11] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[1][11]  ( .G(n17706), .D(n13208), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[1][11] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg2_out_IDEX_reg[11]  ( .D(
        \pipeline/IDEX_Stage/N145 ), .CK(Clk), .Q(n13825), .QN(n17506) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_reg[11]  ( .D(n3868), .CK(Clk), .RN(
        n17704), .Q(n13824), .QN(n7653) );
  DFF_X1 \pipeline/IDEX_Stage/Reg1_out_IDEX_reg[11]  ( .D(
        \pipeline/IDEX_Stage/N113 ), .CK(Clk), .Q(n13823) );
  DFF_X1 \pipeline/MEMWB_Stage/Data_to_RF_reg[9]  ( .D(
        \pipeline/MEMWB_Stage/N20 ), .CK(Clk), .Q(
        \pipeline/data_to_RF_from_WB[9] ), .QN(n17305) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[2][9]  ( .G(n13169), .D(n13202), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[2][9] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[4][9]  ( .G(n13163), .D(n13202), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[4][9] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[6][9]  ( .G(n13157), .D(n13202), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[6][9] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[8][9]  ( .G(n13151), .D(n13202), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[8][9] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[10][9]  ( .G(n13145), .D(n13202), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[10][9] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[12][9]  ( .G(n13139), .D(n13202), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[12][9] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[14][9]  ( .G(n13133), .D(n13202), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[14][9] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[16][9]  ( .G(n13127), .D(n13202), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[16][9] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[18][9]  ( .G(n13121), .D(n13202), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[18][9] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[20][9]  ( .G(n13115), .D(n13202), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[20][9] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[22][9]  ( .G(n13109), .D(n13202), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[22][9] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[24][9]  ( .G(n13103), .D(n13202), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[24][9] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[26][9]  ( .G(n13097), .D(n13202), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[26][9] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[28][9]  ( .G(n13091), .D(n13202), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[28][9] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[30][9]  ( .G(n13085), .D(n13202), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[30][9] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[31][9]  ( .G(n13082), .D(n13202), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[31][9] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[29][9]  ( .G(n13088), .D(n13202), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[29][9] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[27][9]  ( .G(n13094), .D(n13202), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[27][9] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[25][9]  ( .G(n13100), .D(n13202), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[25][9] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[23][9]  ( .G(n13106), .D(n13202), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[23][9] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[21][9]  ( .G(n13112), .D(n13202), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[21][9] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[19][9]  ( .G(n13118), .D(n13202), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[19][9] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[17][9]  ( .G(n13124), .D(n13202), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[17][9] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[15][9]  ( .G(n13130), .D(n13202), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[15][9] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[13][9]  ( .G(n13136), .D(n13202), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[13][9] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[11][9]  ( .G(n13142), .D(n13202), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[11][9] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[9][9]  ( .G(n13148), .D(n13202), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[9][9] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[7][9]  ( .G(n13154), .D(n13202), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[7][9] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[5][9]  ( .G(n13160), .D(n13202), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[5][9] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[3][9]  ( .G(n13166), .D(n13202), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[3][9] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[1][9]  ( .G(n13172), .D(n13202), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[1][9] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg2_out_IDEX_reg[9]  ( .D(
        \pipeline/IDEX_Stage/N143 ), .CK(Clk), .Q(n13822), .QN(n17504) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_reg[9]  ( .D(n3866), .CK(Clk), .RN(
        n17704), .Q(n13821), .QN(n7652) );
  DFF_X1 \pipeline/IDEX_Stage/Reg1_out_IDEX_reg[9]  ( .D(
        \pipeline/IDEX_Stage/N111 ), .CK(Clk), .Q(n13820) );
  DFF_X1 \pipeline/EXMEM_stage/DataToMem_out_EXMEM_reg[9]  ( .D(
        \pipeline/EXMEM_stage/N48 ), .CK(Clk), .Q(n13819) );
  DLH_X1 \DataMem/Mem_reg[7][9]  ( .G(n13079), .D(\DataMem/N2115 ), .Q(
        \DataMem/Mem[7][9] ) );
  DLH_X1 \DataMem/Mem_reg[6][9]  ( .G(n13076), .D(\DataMem/N2051 ), .Q(
        \DataMem/Mem[6][9] ) );
  DLH_X1 \DataMem/Mem_reg[5][9]  ( .G(n13073), .D(\DataMem/N1987 ), .Q(
        \DataMem/Mem[5][9] ) );
  DLH_X1 \DataMem/Mem_reg[4][9]  ( .G(n13070), .D(\DataMem/N1923 ), .Q(
        \DataMem/Mem[4][9] ) );
  DLH_X1 \DataMem/Mem_reg[3][9]  ( .G(n13067), .D(\DataMem/N1859 ), .Q(
        \DataMem/Mem[3][9] ) );
  DLH_X1 \DataMem/Mem_reg[2][9]  ( .G(n13064), .D(\DataMem/N1795 ), .Q(
        \DataMem/Mem[2][9] ) );
  DLH_X1 \DataMem/Mem_reg[1][9]  ( .G(n13061), .D(\DataMem/N1731 ), .Q(
        \DataMem/Mem[1][9] ) );
  DLH_X1 \DataMem/Mem_reg[0][9]  ( .G(n13058), .D(\DataMem/N1667 ), .Q(
        \DataMem/Mem[0][9] ) );
  DLL_X1 \DataMem/Dataout_reg[9]  ( .D(\DataMem/N2188 ), .GN(n13055), .Q(
        \DataMem/N2322 ) );
  DFF_X1 \pipeline/EXMEM_stage/DataToMem_out_EXMEM_reg[11]  ( .D(
        \pipeline/EXMEM_stage/N50 ), .CK(Clk), .Q(n13818) );
  DLH_X1 \DataMem/Mem_reg[7][11]  ( .G(n13079), .D(\DataMem/N2119 ), .Q(
        \DataMem/Mem[7][11] ) );
  DLH_X1 \DataMem/Mem_reg[6][11]  ( .G(n13076), .D(\DataMem/N2055 ), .Q(
        \DataMem/Mem[6][11] ) );
  DLH_X1 \DataMem/Mem_reg[5][11]  ( .G(n13073), .D(\DataMem/N1991 ), .Q(
        \DataMem/Mem[5][11] ) );
  DLH_X1 \DataMem/Mem_reg[4][11]  ( .G(n13070), .D(\DataMem/N1927 ), .Q(
        \DataMem/Mem[4][11] ) );
  DLH_X1 \DataMem/Mem_reg[3][11]  ( .G(n13067), .D(\DataMem/N1863 ), .Q(
        \DataMem/Mem[3][11] ) );
  DLH_X1 \DataMem/Mem_reg[2][11]  ( .G(n13064), .D(\DataMem/N1799 ), .Q(
        \DataMem/Mem[2][11] ) );
  DLH_X1 \DataMem/Mem_reg[1][11]  ( .G(n13061), .D(\DataMem/N1735 ), .Q(
        \DataMem/Mem[1][11] ) );
  DLH_X1 \DataMem/Mem_reg[0][11]  ( .G(n13058), .D(\DataMem/N1671 ), .Q(
        \DataMem/Mem[0][11] ) );
  DLL_X1 \DataMem/Dataout_reg[11]  ( .D(\DataMem/N2194 ), .GN(n13055), .Q(
        \DataMem/N2316 ) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_reg[10]  ( .D(n3864), .CK(Clk), .RN(
        n17705), .Q(n13817), .QN(n7651) );
  DFF_X1 \pipeline/EXMEM_stage/DataToMem_out_EXMEM_reg[10]  ( .D(
        \pipeline/EXMEM_stage/N49 ), .CK(Clk), .Q(n13816) );
  DLH_X1 \DataMem/Mem_reg[7][10]  ( .G(n13079), .D(\DataMem/N2117 ), .Q(
        \DataMem/Mem[7][10] ) );
  DLH_X1 \DataMem/Mem_reg[6][10]  ( .G(n13076), .D(\DataMem/N2053 ), .Q(
        \DataMem/Mem[6][10] ) );
  DLH_X1 \DataMem/Mem_reg[5][10]  ( .G(n13073), .D(\DataMem/N1989 ), .Q(
        \DataMem/Mem[5][10] ) );
  DLH_X1 \DataMem/Mem_reg[4][10]  ( .G(n13070), .D(\DataMem/N1925 ), .Q(
        \DataMem/Mem[4][10] ) );
  DLH_X1 \DataMem/Mem_reg[3][10]  ( .G(n13067), .D(\DataMem/N1861 ), .Q(
        \DataMem/Mem[3][10] ) );
  DLH_X1 \DataMem/Mem_reg[2][10]  ( .G(n13064), .D(\DataMem/N1797 ), .Q(
        \DataMem/Mem[2][10] ) );
  DLH_X1 \DataMem/Mem_reg[1][10]  ( .G(n13061), .D(\DataMem/N1733 ), .Q(
        \DataMem/Mem[1][10] ) );
  DLH_X1 \DataMem/Mem_reg[0][12]  ( .G(n13058), .D(\DataMem/N1673 ), .Q(
        \DataMem/Mem[0][12] ) );
  DLL_X1 \DataMem/Dataout_reg[12]  ( .D(\DataMem/N2197 ), .GN(n13055), .Q(
        \DataMem/N2313 ) );
  DFF_X1 \pipeline/MEMWB_Stage/Data_to_RF_reg[12]  ( .D(
        \pipeline/MEMWB_Stage/N23 ), .CK(Clk), .Q(
        \pipeline/data_to_RF_from_WB[12] ), .QN(n17395) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[2][12]  ( .G(n13169), .D(n13211), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[2][12] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[4][12]  ( .G(n13163), .D(n13211), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[4][12] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[6][12]  ( .G(n13157), .D(n13211), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[6][12] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[8][12]  ( .G(n13151), .D(n13211), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[8][12] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[10][12]  ( .G(n13145), .D(n13211), .Q(\pipeline/RegFile_DEC_WB/RegBank[10][12] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[12][12]  ( .G(n13139), .D(n13211), .Q(\pipeline/RegFile_DEC_WB/RegBank[12][12] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[14][12]  ( .G(n13133), .D(n13211), .Q(\pipeline/RegFile_DEC_WB/RegBank[14][12] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[16][12]  ( .G(n13127), .D(n13211), .Q(\pipeline/RegFile_DEC_WB/RegBank[16][12] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[18][12]  ( .G(n13121), .D(n13211), .Q(\pipeline/RegFile_DEC_WB/RegBank[18][12] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[20][12]  ( .G(n13115), .D(n13211), .Q(\pipeline/RegFile_DEC_WB/RegBank[20][12] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[22][12]  ( .G(n13109), .D(n13211), .Q(\pipeline/RegFile_DEC_WB/RegBank[22][12] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[24][12]  ( .G(n13103), .D(n13211), .Q(\pipeline/RegFile_DEC_WB/RegBank[24][12] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[26][12]  ( .G(n13097), .D(n13211), .Q(\pipeline/RegFile_DEC_WB/RegBank[26][12] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[28][12]  ( .G(n13091), .D(n13211), .Q(\pipeline/RegFile_DEC_WB/RegBank[28][12] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[30][12]  ( .G(n13085), .D(n13211), .Q(\pipeline/RegFile_DEC_WB/RegBank[30][12] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[31][12]  ( .G(n13082), .D(n13211), .Q(\pipeline/RegFile_DEC_WB/RegBank[31][12] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[29][12]  ( .G(n13088), .D(n13211), .Q(\pipeline/RegFile_DEC_WB/RegBank[29][12] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[27][12]  ( .G(n13094), .D(n13211), .Q(\pipeline/RegFile_DEC_WB/RegBank[27][12] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[25][12]  ( .G(n13100), .D(n13211), .Q(\pipeline/RegFile_DEC_WB/RegBank[25][12] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[23][12]  ( .G(n13106), .D(n13211), .Q(\pipeline/RegFile_DEC_WB/RegBank[23][12] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[21][12]  ( .G(n13112), .D(n13211), .Q(\pipeline/RegFile_DEC_WB/RegBank[21][12] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[19][12]  ( .G(n13118), .D(n13211), .Q(\pipeline/RegFile_DEC_WB/RegBank[19][12] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[17][12]  ( .G(n13124), .D(n13211), .Q(\pipeline/RegFile_DEC_WB/RegBank[17][12] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[15][12]  ( .G(n13130), .D(n13211), .Q(\pipeline/RegFile_DEC_WB/RegBank[15][12] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[13][12]  ( .G(n13136), .D(n13211), .Q(\pipeline/RegFile_DEC_WB/RegBank[13][12] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[11][12]  ( .G(n13142), .D(n13211), .Q(\pipeline/RegFile_DEC_WB/RegBank[11][12] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[9][12]  ( .G(n13148), .D(n13211), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[9][12] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[7][12]  ( .G(n13154), .D(n13211), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[7][12] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[5][12]  ( .G(n13160), .D(n13211), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[5][12] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[3][12]  ( .G(n13166), .D(n13211), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[3][12] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[1][12]  ( .G(n13172), .D(n13211), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[1][12] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg2_out_IDEX_reg[12]  ( .D(
        \pipeline/IDEX_Stage/N146 ), .CK(Clk), .Q(n13815), .QN(n17507) );
  DFF_X1 \pipeline/IDEX_Stage/Reg1_out_IDEX_reg[12]  ( .D(
        \pipeline/IDEX_Stage/N114 ), .CK(Clk), .Q(n13814) );
  DFF_X1 \pipeline/EXMEM_stage/ALUres_MEMaddr_out_EXMEM_reg[12]  ( .D(
        \pipeline/EXMEM_stage/N19 ), .CK(Clk), .Q(
        \pipeline/Alu_Out_Addr_to_mem[12] ) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_reg[12]  ( .D(n3862), .CK(Clk), .RN(
        n17705), .Q(n13813), .QN(n7650) );
  DFF_X1 \pipeline/EXMEM_stage/DataToMem_out_EXMEM_reg[12]  ( .D(
        \pipeline/EXMEM_stage/N51 ), .CK(Clk), .Q(n13812) );
  DLH_X1 \DataMem/Mem_reg[7][12]  ( .G(n13079), .D(\DataMem/N2121 ), .Q(
        \DataMem/Mem[7][12] ) );
  DLH_X1 \DataMem/Mem_reg[6][12]  ( .G(n13076), .D(\DataMem/N2057 ), .Q(
        \DataMem/Mem[6][12] ) );
  DLH_X1 \DataMem/Mem_reg[5][12]  ( .G(n13073), .D(\DataMem/N1993 ), .Q(
        \DataMem/Mem[5][12] ) );
  DLH_X1 \DataMem/Mem_reg[4][12]  ( .G(n13070), .D(\DataMem/N1929 ), .Q(
        \DataMem/Mem[4][12] ) );
  DLH_X1 \DataMem/Mem_reg[3][12]  ( .G(n13067), .D(\DataMem/N1865 ), .Q(
        \DataMem/Mem[3][12] ) );
  DLH_X1 \DataMem/Mem_reg[2][12]  ( .G(n13064), .D(\DataMem/N1801 ), .Q(
        \DataMem/Mem[2][12] ) );
  DLH_X1 \DataMem/Mem_reg[1][12]  ( .G(n13061), .D(\DataMem/N1737 ), .Q(
        \DataMem/Mem[1][12] ) );
  DFF_X1 \pipeline/MEMWB_Stage/Data_to_RF_reg[2]  ( .D(
        \pipeline/MEMWB_Stage/N13 ), .CK(Clk), .Q(
        \pipeline/data_to_RF_from_WB[2] ), .QN(n17369) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[2][2]  ( .G(n17707), .D(n13181), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[2][2] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[4][2]  ( .G(n17709), .D(n13181), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[4][2] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[6][2]  ( .G(n17711), .D(n13181), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[6][2] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[8][2]  ( .G(n17713), .D(n13181), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[8][2] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[10][2]  ( .G(n17715), .D(n13181), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[10][2] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[12][2]  ( .G(n17717), .D(n13181), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[12][2] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[14][2]  ( .G(n17719), .D(n13181), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[14][2] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[16][2]  ( .G(n17721), .D(n13181), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[16][2] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[18][2]  ( .G(n17723), .D(n13181), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[18][2] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[20][2]  ( .G(n17725), .D(n13181), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[20][2] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[22][2]  ( .G(n17727), .D(n13181), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[22][2] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[24][2]  ( .G(n17729), .D(n13181), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[24][2] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[26][2]  ( .G(n17731), .D(n13181), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[26][2] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[28][2]  ( .G(n17733), .D(n13181), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[28][2] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[30][2]  ( .G(n17735), .D(n13181), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[30][2] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[31][2]  ( .G(n17736), .D(n13181), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[31][2] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[29][2]  ( .G(n17734), .D(n13181), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[29][2] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[27][2]  ( .G(n17732), .D(n13181), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[27][2] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[25][2]  ( .G(n17730), .D(n13181), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[25][2] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[23][2]  ( .G(n17728), .D(n13181), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[23][2] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[21][2]  ( .G(n17726), .D(n13181), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[21][2] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[19][2]  ( .G(n17724), .D(n13181), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[19][2] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[17][2]  ( .G(n17722), .D(n13181), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[17][2] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[15][2]  ( .G(n17720), .D(n13181), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[15][2] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[13][2]  ( .G(n17718), .D(n13181), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[13][2] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[11][2]  ( .G(n17716), .D(n13181), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[11][2] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[9][2]  ( .G(n17714), .D(n13181), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[9][2] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[7][2]  ( .G(n17712), .D(n13181), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[7][2] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[5][2]  ( .G(n17710), .D(n13181), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[5][2] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[3][2]  ( .G(n17708), .D(n13181), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[3][2] ) );
  DLH_X1 \pipeline/RegFile_DEC_WB/RegBank_reg[1][2]  ( .G(n17706), .D(n13181), 
        .Q(\pipeline/RegFile_DEC_WB/RegBank[1][2] ) );
  DFF_X1 \pipeline/IDEX_Stage/Reg2_out_IDEX_reg[2]  ( .D(
        \pipeline/IDEX_Stage/N136 ), .CK(Clk), .Q(n13811), .QN(n17497) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_reg[2]  ( .D(n3860), .CK(Clk), .RN(
        n17705), .Q(n13810), .QN(n7649) );
  DFF_X1 \pipeline/IDEX_Stage/Reg1_out_IDEX_reg[2]  ( .D(
        \pipeline/IDEX_Stage/N104 ), .CK(Clk), .Q(n13809) );
  DFF_X1 \pipeline/EXMEM_stage/DataToMem_out_EXMEM_reg[2]  ( .D(
        \pipeline/EXMEM_stage/N41 ), .CK(Clk), .Q(n13808) );
  DLH_X1 \DataMem/Mem_reg[7][2]  ( .G(n13079), .D(\DataMem/N2101 ), .Q(
        \DataMem/Mem[7][2] ) );
  DLH_X1 \DataMem/Mem_reg[6][2]  ( .G(n13076), .D(\DataMem/N2037 ), .Q(
        \DataMem/Mem[6][2] ) );
  DLH_X1 \DataMem/Mem_reg[5][2]  ( .G(n13073), .D(\DataMem/N1973 ), .Q(
        \DataMem/Mem[5][2] ) );
  DLH_X1 \DataMem/Mem_reg[4][2]  ( .G(n13070), .D(\DataMem/N1909 ), .Q(
        \DataMem/Mem[4][2] ) );
  DLH_X1 \DataMem/Mem_reg[3][2]  ( .G(n13067), .D(\DataMem/N1845 ), .Q(
        \DataMem/Mem[3][2] ) );
  DLH_X1 \DataMem/Mem_reg[2][2]  ( .G(n13064), .D(\DataMem/N1781 ), .Q(
        \DataMem/Mem[2][2] ) );
  DLH_X1 \DataMem/Mem_reg[1][2]  ( .G(n13061), .D(\DataMem/N1717 ), .Q(
        \DataMem/Mem[1][2] ) );
  DLH_X1 \DataMem/Mem_reg[0][2]  ( .G(n13058), .D(\DataMem/N1653 ), .Q(
        \DataMem/Mem[0][2] ) );
  DLL_X1 \DataMem/Dataout_reg[2]  ( .D(\DataMem/N2167 ), .GN(n17098), .Q(
        \DataMem/N2343 ) );
  DFF_X1 \pipeline/EXMEM_stage/DataToMem_out_EXMEM_reg[3]  ( .D(
        \pipeline/EXMEM_stage/N42 ), .CK(Clk), .Q(n13807) );
  DLH_X1 \DataMem/Mem_reg[7][3]  ( .G(n13079), .D(\DataMem/N2103 ), .Q(
        \DataMem/Mem[7][3] ) );
  DLH_X1 \DataMem/Mem_reg[6][3]  ( .G(n13076), .D(\DataMem/N2039 ), .Q(
        \DataMem/Mem[6][3] ) );
  DLH_X1 \DataMem/Mem_reg[5][3]  ( .G(n13073), .D(\DataMem/N1975 ), .Q(
        \DataMem/Mem[5][3] ) );
  DLH_X1 \DataMem/Mem_reg[4][3]  ( .G(n13070), .D(\DataMem/N1911 ), .Q(
        \DataMem/Mem[4][3] ) );
  DLH_X1 \DataMem/Mem_reg[3][3]  ( .G(n13067), .D(\DataMem/N1847 ), .Q(
        \DataMem/Mem[3][3] ) );
  DLH_X1 \DataMem/Mem_reg[2][3]  ( .G(n13064), .D(\DataMem/N1783 ), .Q(
        \DataMem/Mem[2][3] ) );
  DLH_X1 \DataMem/Mem_reg[1][3]  ( .G(n13061), .D(\DataMem/N1719 ), .Q(
        \DataMem/Mem[1][3] ) );
  DLH_X1 \DataMem/Mem_reg[0][3]  ( .G(n13058), .D(\DataMem/N1655 ), .Q(
        \DataMem/Mem[0][3] ) );
  DLL_X1 \DataMem/Dataout_reg[3]  ( .D(\DataMem/N2170 ), .GN(n17098), .Q(
        \DataMem/N2340 ) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_reg[1]  ( .D(n3858), .CK(Clk), .RN(
        n17705), .Q(n13806), .QN(n7648) );
  DFF_X1 \pipeline/EXMEM_stage/DataToMem_out_EXMEM_reg[1]  ( .D(
        \pipeline/EXMEM_stage/N40 ), .CK(Clk), .Q(n13805) );
  DFF_X1 \pipeline/IDEX_Stage/Reg1_out_IDEX_reg[16]  ( .D(
        \pipeline/IDEX_Stage/N118 ), .CK(Clk), .Q(n13804) );
  DFF_X1 \pipeline/EXMEM_stage/DataToMem_out_EXMEM_reg[16]  ( .D(
        \pipeline/EXMEM_stage/N55 ), .CK(Clk), .Q(n13803) );
  DLH_X1 \DataMem/Mem_reg[7][16]  ( .G(n13079), .D(\DataMem/N2129 ), .Q(
        \DataMem/Mem[7][16] ) );
  DLH_X1 \DataMem/Mem_reg[6][16]  ( .G(n13076), .D(\DataMem/N2065 ), .Q(
        \DataMem/Mem[6][16] ) );
  DLH_X1 \DataMem/Mem_reg[5][16]  ( .G(n13073), .D(\DataMem/N2001 ), .Q(
        \DataMem/Mem[5][16] ) );
  DLH_X1 \DataMem/Mem_reg[4][16]  ( .G(n13070), .D(\DataMem/N1937 ), .Q(
        \DataMem/Mem[4][16] ) );
  DLH_X1 \DataMem/Mem_reg[3][16]  ( .G(n13067), .D(\DataMem/N1873 ), .Q(
        \DataMem/Mem[3][16] ) );
  DLH_X1 \DataMem/Mem_reg[2][16]  ( .G(n13064), .D(\DataMem/N1809 ), .Q(
        \DataMem/Mem[2][16] ) );
  DLH_X1 \DataMem/Mem_reg[1][16]  ( .G(n13061), .D(\DataMem/N1745 ), .Q(
        \DataMem/Mem[1][16] ) );
  DLH_X1 \DataMem/Mem_reg[0][16]  ( .G(n13058), .D(\DataMem/N1681 ), .Q(
        \DataMem/Mem[0][16] ) );
  DLL_X1 \DataMem/Dataout_reg[16]  ( .D(\DataMem/N2209 ), .GN(n13055), .Q(
        \DataMem/N2301 ) );
  DFF_X1 \pipeline/EXMEM_stage/DataToMem_out_EXMEM_reg[17]  ( .D(
        \pipeline/EXMEM_stage/N56 ), .CK(Clk), .Q(n13802) );
  DLH_X1 \DataMem/Mem_reg[7][17]  ( .G(n13079), .D(\DataMem/N2131 ), .Q(
        \DataMem/Mem[7][17] ) );
  DLH_X1 \DataMem/Mem_reg[6][17]  ( .G(n13076), .D(\DataMem/N2067 ), .Q(
        \DataMem/Mem[6][17] ) );
  DLH_X1 \DataMem/Mem_reg[5][17]  ( .G(n13073), .D(\DataMem/N2003 ), .Q(
        \DataMem/Mem[5][17] ) );
  DLH_X1 \DataMem/Mem_reg[4][17]  ( .G(n13070), .D(\DataMem/N1939 ), .Q(
        \DataMem/Mem[4][17] ) );
  DLH_X1 \DataMem/Mem_reg[3][17]  ( .G(n13067), .D(\DataMem/N1875 ), .Q(
        \DataMem/Mem[3][17] ) );
  DLH_X1 \DataMem/Mem_reg[2][17]  ( .G(n13064), .D(\DataMem/N1811 ), .Q(
        \DataMem/Mem[2][17] ) );
  DLH_X1 \DataMem/Mem_reg[1][17]  ( .G(n13061), .D(\DataMem/N1747 ), .Q(
        \DataMem/Mem[1][17] ) );
  DLH_X1 \DataMem/Mem_reg[0][17]  ( .G(n13058), .D(\DataMem/N1683 ), .Q(
        \DataMem/Mem[0][17] ) );
  DLL_X1 \DataMem/Dataout_reg[17]  ( .D(\DataMem/N2212 ), .GN(n13055), .Q(
        \DataMem/N2298 ) );
  DFF_X1 \pipeline/EXMEM_stage/DataToMem_out_EXMEM_reg[18]  ( .D(
        \pipeline/EXMEM_stage/N57 ), .CK(Clk), .Q(n13801) );
  DLH_X1 \DataMem/Mem_reg[7][18]  ( .G(n13079), .D(\DataMem/N2133 ), .Q(
        \DataMem/Mem[7][18] ) );
  DLH_X1 \DataMem/Mem_reg[6][18]  ( .G(n13076), .D(\DataMem/N2069 ), .Q(
        \DataMem/Mem[6][18] ) );
  DLH_X1 \DataMem/Mem_reg[5][18]  ( .G(n13073), .D(\DataMem/N2005 ), .Q(
        \DataMem/Mem[5][18] ) );
  DLH_X1 \DataMem/Mem_reg[4][18]  ( .G(n13070), .D(\DataMem/N1941 ), .Q(
        \DataMem/Mem[4][18] ) );
  DLH_X1 \DataMem/Mem_reg[3][18]  ( .G(n13067), .D(\DataMem/N1877 ), .Q(
        \DataMem/Mem[3][18] ) );
  DLH_X1 \DataMem/Mem_reg[2][18]  ( .G(n13064), .D(\DataMem/N1813 ), .Q(
        \DataMem/Mem[2][18] ) );
  DLH_X1 \DataMem/Mem_reg[1][18]  ( .G(n13061), .D(\DataMem/N1749 ), .Q(
        \DataMem/Mem[1][18] ) );
  DLH_X1 \DataMem/Mem_reg[0][18]  ( .G(n13058), .D(\DataMem/N1685 ), .Q(
        \DataMem/Mem[0][18] ) );
  DLL_X1 \DataMem/Dataout_reg[18]  ( .D(\DataMem/N2215 ), .GN(n17098), .Q(
        \DataMem/N2295 ) );
  DFF_X1 \pipeline/EXMEM_stage/DataToMem_out_EXMEM_reg[19]  ( .D(
        \pipeline/EXMEM_stage/N58 ), .CK(Clk), .Q(n13800) );
  DLH_X1 \DataMem/Mem_reg[7][19]  ( .G(n13079), .D(\DataMem/N2135 ), .Q(
        \DataMem/Mem[7][19] ) );
  DLH_X1 \DataMem/Mem_reg[6][19]  ( .G(n13076), .D(\DataMem/N2071 ), .Q(
        \DataMem/Mem[6][19] ) );
  DLH_X1 \DataMem/Mem_reg[5][19]  ( .G(n13073), .D(\DataMem/N2007 ), .Q(
        \DataMem/Mem[5][19] ) );
  DLH_X1 \DataMem/Mem_reg[4][19]  ( .G(n13070), .D(\DataMem/N1943 ), .Q(
        \DataMem/Mem[4][19] ) );
  DLH_X1 \DataMem/Mem_reg[3][19]  ( .G(n13067), .D(\DataMem/N1879 ), .Q(
        \DataMem/Mem[3][19] ) );
  DLH_X1 \DataMem/Mem_reg[2][19]  ( .G(n13064), .D(\DataMem/N1815 ), .Q(
        \DataMem/Mem[2][19] ) );
  DLH_X1 \DataMem/Mem_reg[1][19]  ( .G(n13061), .D(\DataMem/N1751 ), .Q(
        \DataMem/Mem[1][19] ) );
  DLH_X1 \DataMem/Mem_reg[0][19]  ( .G(n13058), .D(\DataMem/N1687 ), .Q(
        \DataMem/Mem[0][19] ) );
  DLL_X1 \DataMem/Dataout_reg[19]  ( .D(\DataMem/N2218 ), .GN(n13055), .Q(
        \DataMem/N2292 ) );
  DFF_X1 \pipeline/EXMEM_stage/DataToMem_out_EXMEM_reg[20]  ( .D(
        \pipeline/EXMEM_stage/N59 ), .CK(Clk), .Q(n13799) );
  DLH_X1 \DataMem/Mem_reg[7][20]  ( .G(n13079), .D(\DataMem/N2137 ), .Q(
        \DataMem/Mem[7][20] ) );
  DLH_X1 \DataMem/Mem_reg[6][20]  ( .G(n13076), .D(\DataMem/N2073 ), .Q(
        \DataMem/Mem[6][20] ) );
  DLH_X1 \DataMem/Mem_reg[5][20]  ( .G(n13073), .D(\DataMem/N2009 ), .Q(
        \DataMem/Mem[5][20] ) );
  DLH_X1 \DataMem/Mem_reg[4][20]  ( .G(n13070), .D(\DataMem/N1945 ), .Q(
        \DataMem/Mem[4][20] ) );
  DLH_X1 \DataMem/Mem_reg[3][20]  ( .G(n13067), .D(\DataMem/N1881 ), .Q(
        \DataMem/Mem[3][20] ) );
  DLH_X1 \DataMem/Mem_reg[2][20]  ( .G(n13064), .D(\DataMem/N1817 ), .Q(
        \DataMem/Mem[2][20] ) );
  DLH_X1 \DataMem/Mem_reg[1][20]  ( .G(n13061), .D(\DataMem/N1753 ), .Q(
        \DataMem/Mem[1][20] ) );
  DLH_X1 \DataMem/Mem_reg[0][20]  ( .G(n13058), .D(\DataMem/N1689 ), .Q(
        \DataMem/Mem[0][20] ) );
  DLL_X1 \DataMem/Dataout_reg[20]  ( .D(\DataMem/N2221 ), .GN(n17098), .Q(
        \DataMem/N2289 ) );
  DFF_X1 \pipeline/EXMEM_stage/DataToMem_out_EXMEM_reg[21]  ( .D(
        \pipeline/EXMEM_stage/N60 ), .CK(Clk), .Q(n13798) );
  DLH_X1 \DataMem/Mem_reg[7][21]  ( .G(n13079), .D(\DataMem/N2139 ), .Q(
        \DataMem/Mem[7][21] ) );
  DLH_X1 \DataMem/Mem_reg[6][21]  ( .G(n13076), .D(\DataMem/N2075 ), .Q(
        \DataMem/Mem[6][21] ) );
  DLH_X1 \DataMem/Mem_reg[5][21]  ( .G(n13073), .D(\DataMem/N2011 ), .Q(
        \DataMem/Mem[5][21] ) );
  DLH_X1 \DataMem/Mem_reg[4][21]  ( .G(n13070), .D(\DataMem/N1947 ), .Q(
        \DataMem/Mem[4][21] ) );
  DLH_X1 \DataMem/Mem_reg[3][21]  ( .G(n13067), .D(\DataMem/N1883 ), .Q(
        \DataMem/Mem[3][21] ) );
  DLH_X1 \DataMem/Mem_reg[2][21]  ( .G(n13064), .D(\DataMem/N1819 ), .Q(
        \DataMem/Mem[2][21] ) );
  DLH_X1 \DataMem/Mem_reg[1][21]  ( .G(n13061), .D(\DataMem/N1755 ), .Q(
        \DataMem/Mem[1][21] ) );
  DLH_X1 \DataMem/Mem_reg[0][21]  ( .G(n13058), .D(\DataMem/N1691 ), .Q(
        \DataMem/Mem[0][21] ) );
  DLL_X1 \DataMem/Dataout_reg[21]  ( .D(\DataMem/N2224 ), .GN(n17098), .Q(
        \DataMem/N2286 ) );
  DFF_X1 \pipeline/EXMEM_stage/DataToMem_out_EXMEM_reg[22]  ( .D(
        \pipeline/EXMEM_stage/N61 ), .CK(Clk), .Q(n13797) );
  DLH_X1 \DataMem/Mem_reg[7][22]  ( .G(n13079), .D(\DataMem/N2141 ), .Q(
        \DataMem/Mem[7][22] ) );
  DLH_X1 \DataMem/Mem_reg[6][22]  ( .G(n13076), .D(\DataMem/N2077 ), .Q(
        \DataMem/Mem[6][22] ) );
  DLH_X1 \DataMem/Mem_reg[5][22]  ( .G(n13073), .D(\DataMem/N2013 ), .Q(
        \DataMem/Mem[5][22] ) );
  DLH_X1 \DataMem/Mem_reg[4][22]  ( .G(n13070), .D(\DataMem/N1949 ), .Q(
        \DataMem/Mem[4][22] ) );
  DLH_X1 \DataMem/Mem_reg[3][22]  ( .G(n13067), .D(\DataMem/N1885 ), .Q(
        \DataMem/Mem[3][22] ) );
  DLH_X1 \DataMem/Mem_reg[2][22]  ( .G(n13064), .D(\DataMem/N1821 ), .Q(
        \DataMem/Mem[2][22] ) );
  DLH_X1 \DataMem/Mem_reg[1][22]  ( .G(n13061), .D(\DataMem/N1757 ), .Q(
        \DataMem/Mem[1][22] ) );
  DLH_X1 \DataMem/Mem_reg[0][22]  ( .G(n13058), .D(\DataMem/N1693 ), .Q(
        \DataMem/Mem[0][22] ) );
  DLL_X1 \DataMem/Dataout_reg[22]  ( .D(\DataMem/N2227 ), .GN(n13055), .Q(
        \DataMem/N2283 ) );
  DFF_X1 \pipeline/EXMEM_stage/DataToMem_out_EXMEM_reg[23]  ( .D(
        \pipeline/EXMEM_stage/N62 ), .CK(Clk), .Q(n13796) );
  DLH_X1 \DataMem/Mem_reg[7][23]  ( .G(n13079), .D(\DataMem/N2143 ), .Q(
        \DataMem/Mem[7][23] ) );
  DLH_X1 \DataMem/Mem_reg[6][23]  ( .G(n13076), .D(\DataMem/N2079 ), .Q(
        \DataMem/Mem[6][23] ) );
  DLH_X1 \DataMem/Mem_reg[5][23]  ( .G(n13073), .D(\DataMem/N2015 ), .Q(
        \DataMem/Mem[5][23] ) );
  DLH_X1 \DataMem/Mem_reg[4][23]  ( .G(n13070), .D(\DataMem/N1951 ), .Q(
        \DataMem/Mem[4][23] ) );
  DLH_X1 \DataMem/Mem_reg[3][23]  ( .G(n13067), .D(\DataMem/N1887 ), .Q(
        \DataMem/Mem[3][23] ) );
  DLH_X1 \DataMem/Mem_reg[2][23]  ( .G(n13064), .D(\DataMem/N1823 ), .Q(
        \DataMem/Mem[2][23] ) );
  DLH_X1 \DataMem/Mem_reg[1][23]  ( .G(n13061), .D(\DataMem/N1759 ), .Q(
        \DataMem/Mem[1][23] ) );
  DLH_X1 \DataMem/Mem_reg[0][23]  ( .G(n13058), .D(\DataMem/N1695 ), .Q(
        \DataMem/Mem[0][23] ) );
  DLL_X1 \DataMem/Dataout_reg[23]  ( .D(\DataMem/N2230 ), .GN(n13055), .Q(
        \DataMem/N2280 ) );
  DFF_X1 \pipeline/EXMEM_stage/DataToMem_out_EXMEM_reg[25]  ( .D(
        \pipeline/EXMEM_stage/N64 ), .CK(Clk), .Q(n13795) );
  DLH_X1 \DataMem/Mem_reg[7][25]  ( .G(n13079), .D(\DataMem/N2147 ), .Q(
        \DataMem/Mem[7][25] ) );
  DLH_X1 \DataMem/Mem_reg[6][25]  ( .G(n13076), .D(\DataMem/N2083 ), .Q(
        \DataMem/Mem[6][25] ) );
  DLH_X1 \DataMem/Mem_reg[5][25]  ( .G(n13073), .D(\DataMem/N2019 ), .Q(
        \DataMem/Mem[5][25] ) );
  DLH_X1 \DataMem/Mem_reg[4][25]  ( .G(n13070), .D(\DataMem/N1955 ), .Q(
        \DataMem/Mem[4][25] ) );
  DLH_X1 \DataMem/Mem_reg[3][25]  ( .G(n13067), .D(\DataMem/N1891 ), .Q(
        \DataMem/Mem[3][25] ) );
  DLH_X1 \DataMem/Mem_reg[2][25]  ( .G(n13064), .D(\DataMem/N1827 ), .Q(
        \DataMem/Mem[2][25] ) );
  DLH_X1 \DataMem/Mem_reg[1][25]  ( .G(n13061), .D(\DataMem/N1763 ), .Q(
        \DataMem/Mem[1][25] ) );
  DLH_X1 \DataMem/Mem_reg[0][25]  ( .G(n13058), .D(\DataMem/N1699 ), .Q(
        \DataMem/Mem[0][25] ) );
  DLL_X1 \DataMem/Dataout_reg[25]  ( .D(\DataMem/N2236 ), .GN(n17098), .Q(
        \DataMem/N2274 ) );
  DFF_X1 \pipeline/EXMEM_stage/DataToMem_out_EXMEM_reg[26]  ( .D(
        \pipeline/EXMEM_stage/N65 ), .CK(Clk), .Q(n13794) );
  DLH_X1 \DataMem/Mem_reg[7][26]  ( .G(n13079), .D(\DataMem/N2149 ), .Q(
        \DataMem/Mem[7][26] ) );
  DLH_X1 \DataMem/Mem_reg[6][26]  ( .G(n13076), .D(\DataMem/N2085 ), .Q(
        \DataMem/Mem[6][26] ) );
  DLH_X1 \DataMem/Mem_reg[5][26]  ( .G(n13073), .D(\DataMem/N2021 ), .Q(
        \DataMem/Mem[5][26] ) );
  DLH_X1 \DataMem/Mem_reg[4][26]  ( .G(n13070), .D(\DataMem/N1957 ), .Q(
        \DataMem/Mem[4][26] ) );
  DLH_X1 \DataMem/Mem_reg[3][26]  ( .G(n13067), .D(\DataMem/N1893 ), .Q(
        \DataMem/Mem[3][26] ) );
  DLH_X1 \DataMem/Mem_reg[2][26]  ( .G(n13064), .D(\DataMem/N1829 ), .Q(
        \DataMem/Mem[2][26] ) );
  DLH_X1 \DataMem/Mem_reg[1][26]  ( .G(n13061), .D(\DataMem/N1765 ), .Q(
        \DataMem/Mem[1][26] ) );
  DLH_X1 \DataMem/Mem_reg[0][26]  ( .G(n13058), .D(\DataMem/N1701 ), .Q(
        \DataMem/Mem[0][26] ) );
  DLL_X1 \DataMem/Dataout_reg[26]  ( .D(\DataMem/N2239 ), .GN(n17098), .Q(
        \DataMem/N2271 ) );
  DFF_X1 \pipeline/EXMEM_stage/DataToMem_out_EXMEM_reg[27]  ( .D(
        \pipeline/EXMEM_stage/N66 ), .CK(Clk), .Q(n13793) );
  DLH_X1 \DataMem/Mem_reg[7][27]  ( .G(n13079), .D(\DataMem/N2151 ), .Q(
        \DataMem/Mem[7][27] ) );
  DLH_X1 \DataMem/Mem_reg[6][27]  ( .G(n13076), .D(\DataMem/N2087 ), .Q(
        \DataMem/Mem[6][27] ) );
  DLH_X1 \DataMem/Mem_reg[5][27]  ( .G(n13073), .D(\DataMem/N2023 ), .Q(
        \DataMem/Mem[5][27] ) );
  DLH_X1 \DataMem/Mem_reg[4][27]  ( .G(n13070), .D(\DataMem/N1959 ), .Q(
        \DataMem/Mem[4][27] ) );
  DLH_X1 \DataMem/Mem_reg[3][27]  ( .G(n13067), .D(\DataMem/N1895 ), .Q(
        \DataMem/Mem[3][27] ) );
  DLH_X1 \DataMem/Mem_reg[2][27]  ( .G(n13064), .D(\DataMem/N1831 ), .Q(
        \DataMem/Mem[2][27] ) );
  DLH_X1 \DataMem/Mem_reg[1][27]  ( .G(n13061), .D(\DataMem/N1767 ), .Q(
        \DataMem/Mem[1][27] ) );
  DLH_X1 \DataMem/Mem_reg[0][27]  ( .G(n13058), .D(\DataMem/N1703 ), .Q(
        \DataMem/Mem[0][27] ) );
  DLL_X1 \DataMem/Dataout_reg[27]  ( .D(\DataMem/N2242 ), .GN(n17098), .Q(
        \DataMem/N2268 ) );
  DFF_X1 \pipeline/EXMEM_stage/DataToMem_out_EXMEM_reg[29]  ( .D(
        \pipeline/EXMEM_stage/N68 ), .CK(Clk), .Q(n13792) );
  DLH_X1 \DataMem/Mem_reg[7][29]  ( .G(n13079), .D(\DataMem/N2155 ), .Q(
        \DataMem/Mem[7][29] ) );
  DLH_X1 \DataMem/Mem_reg[6][29]  ( .G(n13076), .D(\DataMem/N2091 ), .Q(
        \DataMem/Mem[6][29] ) );
  DLH_X1 \DataMem/Mem_reg[5][29]  ( .G(n13073), .D(\DataMem/N2027 ), .Q(
        \DataMem/Mem[5][29] ) );
  DLH_X1 \DataMem/Mem_reg[4][29]  ( .G(n13070), .D(\DataMem/N1963 ), .Q(
        \DataMem/Mem[4][29] ) );
  DLH_X1 \DataMem/Mem_reg[3][29]  ( .G(n13067), .D(\DataMem/N1899 ), .Q(
        \DataMem/Mem[3][29] ) );
  DLH_X1 \DataMem/Mem_reg[2][29]  ( .G(n13064), .D(\DataMem/N1835 ), .Q(
        \DataMem/Mem[2][29] ) );
  DLH_X1 \DataMem/Mem_reg[1][29]  ( .G(n13061), .D(\DataMem/N1771 ), .Q(
        \DataMem/Mem[1][29] ) );
  DLH_X1 \DataMem/Mem_reg[0][29]  ( .G(n13058), .D(\DataMem/N1707 ), .Q(
        \DataMem/Mem[0][29] ) );
  DLL_X1 \DataMem/Dataout_reg[29]  ( .D(\DataMem/N2248 ), .GN(n17098), .Q(
        \DataMem/N2262 ) );
  DFF_X1 \pipeline/EXMEM_stage/DataToMem_out_EXMEM_reg[30]  ( .D(
        \pipeline/EXMEM_stage/N69 ), .CK(Clk), .Q(n13791) );
  DLH_X1 \DataMem/Mem_reg[7][30]  ( .G(n13079), .D(\DataMem/N2157 ), .Q(
        \DataMem/Mem[7][30] ) );
  DLH_X1 \DataMem/Mem_reg[6][30]  ( .G(n13076), .D(\DataMem/N2093 ), .Q(
        \DataMem/Mem[6][30] ) );
  DLH_X1 \DataMem/Mem_reg[5][30]  ( .G(n13073), .D(\DataMem/N2029 ), .Q(
        \DataMem/Mem[5][30] ) );
  DLH_X1 \DataMem/Mem_reg[4][30]  ( .G(n13070), .D(\DataMem/N1965 ), .Q(
        \DataMem/Mem[4][30] ) );
  DLH_X1 \DataMem/Mem_reg[3][30]  ( .G(n13067), .D(\DataMem/N1901 ), .Q(
        \DataMem/Mem[3][30] ) );
  DLH_X1 \DataMem/Mem_reg[2][30]  ( .G(n13064), .D(\DataMem/N1837 ), .Q(
        \DataMem/Mem[2][30] ) );
  DLH_X1 \DataMem/Mem_reg[1][30]  ( .G(n13061), .D(\DataMem/N1773 ), .Q(
        \DataMem/Mem[1][30] ) );
  DLH_X1 \DataMem/Mem_reg[0][30]  ( .G(n13058), .D(\DataMem/N1709 ), .Q(
        \DataMem/Mem[0][30] ) );
  DLL_X1 \DataMem/Dataout_reg[30]  ( .D(\DataMem/N2251 ), .GN(n17098), .Q(
        \DataMem/N2259 ) );
  DFF_X1 \pipeline/EXMEM_stage/DataToMem_out_EXMEM_reg[13]  ( .D(
        \pipeline/EXMEM_stage/N52 ), .CK(Clk), .Q(n13790) );
  DLH_X1 \DataMem/Mem_reg[7][13]  ( .G(n13079), .D(\DataMem/N2123 ), .Q(
        \DataMem/Mem[7][13] ) );
  DLH_X1 \DataMem/Mem_reg[6][13]  ( .G(n13076), .D(\DataMem/N2059 ), .Q(
        \DataMem/Mem[6][13] ) );
  DLH_X1 \DataMem/Mem_reg[5][13]  ( .G(n13073), .D(\DataMem/N1995 ), .Q(
        \DataMem/Mem[5][13] ) );
  DLH_X1 \DataMem/Mem_reg[4][13]  ( .G(n13070), .D(\DataMem/N1931 ), .Q(
        \DataMem/Mem[4][13] ) );
  DLH_X1 \DataMem/Mem_reg[3][13]  ( .G(n13067), .D(\DataMem/N1867 ), .Q(
        \DataMem/Mem[3][13] ) );
  DLH_X1 \DataMem/Mem_reg[2][13]  ( .G(n13064), .D(\DataMem/N1803 ), .Q(
        \DataMem/Mem[2][13] ) );
  DLH_X1 \DataMem/Mem_reg[1][13]  ( .G(n13061), .D(\DataMem/N1739 ), .Q(
        \DataMem/Mem[1][13] ) );
  DLH_X1 \DataMem/Mem_reg[0][13]  ( .G(n13058), .D(\DataMem/N1675 ), .Q(
        \DataMem/Mem[0][13] ) );
  DLL_X1 \DataMem/Dataout_reg[13]  ( .D(\DataMem/N2200 ), .GN(n13055), .Q(
        \DataMem/N2310 ) );
  DFF_X1 \pipeline/EXMEM_stage/DataToMem_out_EXMEM_reg[15]  ( .D(
        \pipeline/EXMEM_stage/N54 ), .CK(Clk), .Q(n13789) );
  DLH_X1 \DataMem/Mem_reg[7][15]  ( .G(n13079), .D(\DataMem/N2127 ), .Q(
        \DataMem/Mem[7][15] ) );
  DLH_X1 \DataMem/Mem_reg[6][15]  ( .G(n13076), .D(\DataMem/N2063 ), .Q(
        \DataMem/Mem[6][15] ) );
  DLH_X1 \DataMem/Mem_reg[5][15]  ( .G(n13073), .D(\DataMem/N1999 ), .Q(
        \DataMem/Mem[5][15] ) );
  DLH_X1 \DataMem/Mem_reg[4][15]  ( .G(n13070), .D(\DataMem/N1935 ), .Q(
        \DataMem/Mem[4][15] ) );
  DLH_X1 \DataMem/Mem_reg[3][15]  ( .G(n13067), .D(\DataMem/N1871 ), .Q(
        \DataMem/Mem[3][15] ) );
  DLH_X1 \DataMem/Mem_reg[2][15]  ( .G(n13064), .D(\DataMem/N1807 ), .Q(
        \DataMem/Mem[2][15] ) );
  DLH_X1 \DataMem/Mem_reg[1][15]  ( .G(n13061), .D(\DataMem/N1743 ), .Q(
        \DataMem/Mem[1][15] ) );
  DLH_X1 \DataMem/Mem_reg[0][15]  ( .G(n13058), .D(\DataMem/N1679 ), .Q(
        \DataMem/Mem[0][15] ) );
  DLL_X1 \DataMem/Dataout_reg[15]  ( .D(\DataMem/N2206 ), .GN(n13055), .Q(
        \DataMem/N2304 ) );
  DFF_X1 \pipeline/EXMEM_stage/DataToMem_out_EXMEM_reg[14]  ( .D(
        \pipeline/EXMEM_stage/N53 ), .CK(Clk), .Q(n13788) );
  DLH_X1 \DataMem/Mem_reg[7][14]  ( .G(n13079), .D(\DataMem/N2125 ), .Q(
        \DataMem/Mem[7][14] ) );
  DLH_X1 \DataMem/Mem_reg[6][14]  ( .G(n13076), .D(\DataMem/N2061 ), .Q(
        \DataMem/Mem[6][14] ) );
  DLH_X1 \DataMem/Mem_reg[5][14]  ( .G(n13073), .D(\DataMem/N1997 ), .Q(
        \DataMem/Mem[5][14] ) );
  DLH_X1 \DataMem/Mem_reg[4][14]  ( .G(n13070), .D(\DataMem/N1933 ), .Q(
        \DataMem/Mem[4][14] ) );
  DLH_X1 \DataMem/Mem_reg[3][14]  ( .G(n13067), .D(\DataMem/N1869 ), .Q(
        \DataMem/Mem[3][14] ) );
  DLH_X1 \DataMem/Mem_reg[2][14]  ( .G(n13064), .D(\DataMem/N1805 ), .Q(
        \DataMem/Mem[2][14] ) );
  DLH_X1 \DataMem/Mem_reg[1][14]  ( .G(n13061), .D(\DataMem/N1741 ), .Q(
        \DataMem/Mem[1][14] ) );
  DLH_X1 \DataMem/Mem_reg[0][14]  ( .G(n13058), .D(\DataMem/N1677 ), .Q(
        \DataMem/Mem[0][14] ) );
  DLL_X1 \DataMem/Dataout_reg[14]  ( .D(\DataMem/N2203 ), .GN(n13055), .Q(
        \DataMem/N2307 ) );
  DFF_X1 \pipeline/EXMEM_stage/DataToMem_out_EXMEM_reg[28]  ( .D(
        \pipeline/EXMEM_stage/N67 ), .CK(Clk), .Q(n13787) );
  DLH_X1 \DataMem/Mem_reg[7][28]  ( .G(n13079), .D(\DataMem/N2153 ), .Q(
        \DataMem/Mem[7][28] ) );
  DLH_X1 \DataMem/Mem_reg[6][28]  ( .G(n13076), .D(\DataMem/N2089 ), .Q(
        \DataMem/Mem[6][28] ) );
  DLH_X1 \DataMem/Mem_reg[5][28]  ( .G(n13073), .D(\DataMem/N2025 ), .Q(
        \DataMem/Mem[5][28] ) );
  DLH_X1 \DataMem/Mem_reg[4][28]  ( .G(n13070), .D(\DataMem/N1961 ), .Q(
        \DataMem/Mem[4][28] ) );
  DLH_X1 \DataMem/Mem_reg[3][28]  ( .G(n13067), .D(\DataMem/N1897 ), .Q(
        \DataMem/Mem[3][28] ) );
  DLH_X1 \DataMem/Mem_reg[2][28]  ( .G(n13064), .D(\DataMem/N1833 ), .Q(
        \DataMem/Mem[2][28] ) );
  DLH_X1 \DataMem/Mem_reg[1][28]  ( .G(n13061), .D(\DataMem/N1769 ), .Q(
        \DataMem/Mem[1][28] ) );
  DLH_X1 \DataMem/Mem_reg[0][28]  ( .G(n13058), .D(\DataMem/N1705 ), .Q(
        \DataMem/Mem[0][28] ) );
  DLL_X1 \DataMem/Dataout_reg[28]  ( .D(\DataMem/N2245 ), .GN(n17098), .Q(
        \DataMem/N2265 ) );
  DFF_X1 \pipeline/EXMEM_stage/DataToMem_out_EXMEM_reg[24]  ( .D(
        \pipeline/EXMEM_stage/N63 ), .CK(Clk), .Q(n13786) );
  DLH_X1 \DataMem/Mem_reg[7][24]  ( .G(n13079), .D(\DataMem/N2145 ), .Q(
        \DataMem/Mem[7][24] ) );
  DLH_X1 \DataMem/Mem_reg[6][24]  ( .G(n13076), .D(\DataMem/N2081 ), .Q(
        \DataMem/Mem[6][24] ) );
  DLH_X1 \DataMem/Mem_reg[5][24]  ( .G(n13073), .D(\DataMem/N2017 ), .Q(
        \DataMem/Mem[5][24] ) );
  DLH_X1 \DataMem/Mem_reg[4][24]  ( .G(n13070), .D(\DataMem/N1953 ), .Q(
        \DataMem/Mem[4][24] ) );
  DLH_X1 \DataMem/Mem_reg[3][24]  ( .G(n13067), .D(\DataMem/N1889 ), .Q(
        \DataMem/Mem[3][24] ) );
  DLH_X1 \DataMem/Mem_reg[2][24]  ( .G(n13064), .D(\DataMem/N1825 ), .Q(
        \DataMem/Mem[2][24] ) );
  DLH_X1 \DataMem/Mem_reg[1][24]  ( .G(n13061), .D(\DataMem/N1761 ), .Q(
        \DataMem/Mem[1][24] ) );
  DLH_X1 \DataMem/Mem_reg[0][24]  ( .G(n13058), .D(\DataMem/N1697 ), .Q(
        \DataMem/Mem[0][24] ) );
  DLL_X1 \DataMem/Dataout_reg[24]  ( .D(\DataMem/N2233 ), .GN(n13055), .Q(
        \DataMem/N2277 ) );
  DFF_X1 \pipeline/EXMEM_stage/DataToMem_out_EXMEM_reg[8]  ( .D(
        \pipeline/EXMEM_stage/N47 ), .CK(Clk), .Q(n13785) );
  DLH_X1 \DataMem/Mem_reg[7][8]  ( .G(n13079), .D(\DataMem/N2113 ), .Q(
        \DataMem/Mem[7][8] ) );
  DLH_X1 \DataMem/Mem_reg[6][8]  ( .G(n13076), .D(\DataMem/N2049 ), .Q(
        \DataMem/Mem[6][8] ) );
  DLH_X1 \DataMem/Mem_reg[5][8]  ( .G(n13073), .D(\DataMem/N1985 ), .Q(
        \DataMem/Mem[5][8] ) );
  DLH_X1 \DataMem/Mem_reg[4][8]  ( .G(n13070), .D(\DataMem/N1921 ), .Q(
        \DataMem/Mem[4][8] ) );
  DLH_X1 \DataMem/Mem_reg[3][8]  ( .G(n13067), .D(\DataMem/N1857 ), .Q(
        \DataMem/Mem[3][8] ) );
  DLH_X1 \DataMem/Mem_reg[2][8]  ( .G(n13064), .D(\DataMem/N1793 ), .Q(
        \DataMem/Mem[2][8] ) );
  DLH_X1 \DataMem/Mem_reg[1][8]  ( .G(n13061), .D(\DataMem/N1729 ), .Q(
        \DataMem/Mem[1][8] ) );
  DLH_X1 \DataMem/Mem_reg[0][8]  ( .G(n13058), .D(\DataMem/N1665 ), .Q(
        \DataMem/Mem[0][8] ) );
  DLL_X1 \DataMem/Dataout_reg[8]  ( .D(\DataMem/N2185 ), .GN(n17098), .Q(
        \DataMem/N2325 ) );
  DFF_X1 \pipeline/EXMEM_stage/DataToMem_out_EXMEM_reg[0]  ( .D(
        \pipeline/EXMEM_stage/N39 ), .CK(Clk), .Q(n13784) );
  DLH_X1 \DataMem/Mem_reg[7][0]  ( .G(n13079), .D(\DataMem/N2097 ), .Q(
        \DataMem/Mem[7][0] ) );
  DLH_X1 \DataMem/Mem_reg[6][0]  ( .G(n13076), .D(\DataMem/N2033 ), .Q(
        \DataMem/Mem[6][0] ) );
  DLH_X1 \DataMem/Mem_reg[5][0]  ( .G(n13073), .D(\DataMem/N1969 ), .Q(
        \DataMem/Mem[5][0] ) );
  DLH_X1 \DataMem/Mem_reg[4][0]  ( .G(n13070), .D(\DataMem/N1905 ), .Q(
        \DataMem/Mem[4][0] ) );
  DLH_X1 \DataMem/Mem_reg[3][0]  ( .G(n13067), .D(\DataMem/N1841 ), .Q(
        \DataMem/Mem[3][0] ) );
  DLH_X1 \DataMem/Mem_reg[2][0]  ( .G(n13064), .D(\DataMem/N1777 ), .Q(
        \DataMem/Mem[2][0] ) );
  DLH_X1 \DataMem/Mem_reg[1][0]  ( .G(n13061), .D(\DataMem/N1713 ), .Q(
        \DataMem/Mem[1][0] ) );
  DLH_X1 \DataMem/Mem_reg[0][0]  ( .G(n13058), .D(\DataMem/N1649 ), .Q(
        \DataMem/Mem[0][0] ) );
  DLL_X1 \DataMem/Dataout_reg[0]  ( .D(\DataMem/N2161 ), .GN(n17098), .Q(
        \DataMem/N2349 ) );
  DFF_X1 \pipeline/EXMEM_stage/DataToMem_out_EXMEM_reg[31]  ( .D(
        \pipeline/EXMEM_stage/N70 ), .CK(Clk), .Q(n13783) );
  DLH_X1 \DataMem/Mem_reg[6][31]  ( .G(n13076), .D(\DataMem/N2095 ), .Q(
        \DataMem/Mem[6][31] ) );
  DLH_X1 \DataMem/Mem_reg[5][31]  ( .G(n13073), .D(\DataMem/N2031 ), .Q(
        \DataMem/Mem[5][31] ) );
  DLH_X1 \DataMem/Mem_reg[4][31]  ( .G(n13070), .D(\DataMem/N1967 ), .Q(
        \DataMem/Mem[4][31] ) );
  DLH_X1 \DataMem/Mem_reg[3][31]  ( .G(n13067), .D(\DataMem/N1903 ), .Q(
        \DataMem/Mem[3][31] ) );
  DLH_X1 \DataMem/Mem_reg[2][31]  ( .G(n13064), .D(\DataMem/N1839 ), .Q(
        \DataMem/Mem[2][31] ) );
  DLH_X1 \DataMem/Mem_reg[1][31]  ( .G(n13061), .D(\DataMem/N1775 ), .Q(
        \DataMem/Mem[1][31] ) );
  DLH_X1 \DataMem/Mem_reg[0][31]  ( .G(n13058), .D(\DataMem/N1711 ), .Q(
        \DataMem/Mem[0][31] ) );
  DLL_X1 \pipeline/stageM/Addr_to_Dram_reg[4]  ( .D(
        \pipeline/Alu_Out_Addr_to_mem[4] ), .GN(n12766), .Q(addr_to_dataRam[4]) );
  DFF_X2 \pipeline/IDEX_Stage/EXE_controls_out_IDEX_reg[1]  ( .D(
        \pipeline/IDEX_Stage/N94 ), .CK(Clk), .Q(
        \pipeline/stageE/EXE_ALU/add_alu/sCout[0] ), .QN(n17381) );
  DLL_X1 \pipeline/stageM/Addr_to_Dram_reg[3]  ( .D(
        \pipeline/Alu_Out_Addr_to_mem[3] ), .GN(n17155), .Q(addr_to_dataRam[3]) );
  DLL_X1 \pipeline/stageM/Addr_to_Dram_reg[2]  ( .D(
        \pipeline/Alu_Out_Addr_to_mem[2] ), .GN(n12766), .Q(addr_to_dataRam[2]) );
  TINV_X1 U4372 ( .I(n7676), .EN(\pipeline/stageF/PC_reg/N0 ), .ZN(
        addr_to_iram[31]) );
  TINV_X1 U4374 ( .I(n7649), .EN(\pipeline/stageF/PC_reg/N29 ), .ZN(
        addr_to_iram[2]) );
  TINV_X1 U4375 ( .I(n7659), .EN(\pipeline/stageF/PC_reg/N31 ), .ZN(
        \pipeline/stageF/PC_plus4/N7 ) );
  TINV_X1 U4376 ( .I(n7648), .EN(\pipeline/stageF/PC_reg/N30 ), .ZN(
        \pipeline/stageF/PC_plus4/N8 ) );
  TINV_X1 U4377 ( .I(n7658), .EN(\pipeline/stageF/PC_reg/N28 ), .ZN(
        addr_to_iram[3]) );
  TINV_X1 U4378 ( .I(n7656), .EN(\pipeline/stageF/PC_reg/N27 ), .ZN(
        addr_to_iram[4]) );
  TINV_X1 U4379 ( .I(n7655), .EN(\pipeline/stageF/PC_reg/N26 ), .ZN(
        addr_to_iram[5]) );
  TINV_X1 U4380 ( .I(n7654), .EN(\pipeline/stageF/PC_reg/N25 ), .ZN(
        addr_to_iram[6]) );
  TINV_X1 U4381 ( .I(n7657), .EN(\pipeline/stageF/PC_reg/N24 ), .ZN(
        addr_to_iram[7]) );
  TINV_X1 U4382 ( .I(n7660), .EN(\pipeline/stageF/PC_reg/N23 ), .ZN(
        addr_to_iram[8]) );
  TINV_X1 U4383 ( .I(n7652), .EN(\pipeline/stageF/PC_reg/N22 ), .ZN(
        addr_to_iram[9]) );
  TINV_X1 U4384 ( .I(n7651), .EN(\pipeline/stageF/PC_reg/N21 ), .ZN(
        addr_to_iram[10]) );
  TINV_X1 U4385 ( .I(n7653), .EN(\pipeline/stageF/PC_reg/N20 ), .ZN(
        addr_to_iram[11]) );
  TINV_X1 U4386 ( .I(n7650), .EN(\pipeline/stageF/PC_reg/N19 ), .ZN(
        addr_to_iram[12]) );
  TINV_X1 U4387 ( .I(n7661), .EN(\pipeline/stageF/PC_reg/N18 ), .ZN(
        addr_to_iram[13]) );
  TINV_X1 U4388 ( .I(n7662), .EN(\pipeline/stageF/PC_reg/N17 ), .ZN(
        addr_to_iram[14]) );
  TINV_X1 U4389 ( .I(n7663), .EN(\pipeline/stageF/PC_reg/N16 ), .ZN(
        addr_to_iram[15]) );
  TINV_X1 U4390 ( .I(n7711), .EN(\pipeline/stageF/PC_reg/N15 ), .ZN(
        addr_to_iram[16]) );
  TINV_X1 U4391 ( .I(n7664), .EN(\pipeline/stageF/PC_reg/N14 ), .ZN(
        addr_to_iram[17]) );
  TINV_X1 U4392 ( .I(n7665), .EN(\pipeline/stageF/PC_reg/N13 ), .ZN(
        addr_to_iram[18]) );
  TINV_X1 U4393 ( .I(n7666), .EN(\pipeline/stageF/PC_reg/N12 ), .ZN(
        addr_to_iram[19]) );
  TINV_X1 U4394 ( .I(n7667), .EN(\pipeline/stageF/PC_reg/N11 ), .ZN(
        addr_to_iram[20]) );
  TINV_X1 U4395 ( .I(n7668), .EN(\pipeline/stageF/PC_reg/N10 ), .ZN(
        addr_to_iram[21]) );
  TINV_X1 U4396 ( .I(n7669), .EN(\pipeline/stageF/PC_reg/N9 ), .ZN(
        addr_to_iram[22]) );
  TINV_X1 U4397 ( .I(n7670), .EN(\pipeline/stageF/PC_reg/N8 ), .ZN(
        addr_to_iram[23]) );
  TINV_X1 U4398 ( .I(n7671), .EN(\pipeline/stageF/PC_reg/N7 ), .ZN(
        addr_to_iram[24]) );
  TINV_X1 U4399 ( .I(n7672), .EN(\pipeline/stageF/PC_reg/N6 ), .ZN(
        addr_to_iram[25]) );
  TINV_X1 U4400 ( .I(n7673), .EN(\pipeline/stageF/PC_reg/N5 ), .ZN(
        addr_to_iram[26]) );
  TINV_X1 U4401 ( .I(n7674), .EN(\pipeline/stageF/PC_reg/N4 ), .ZN(
        addr_to_iram[27]) );
  TINV_X1 U4402 ( .I(n7675), .EN(\pipeline/stageF/PC_reg/N3 ), .ZN(
        addr_to_iram[28]) );
  TINV_X1 U4403 ( .I(n7709), .EN(\pipeline/stageF/PC_reg/N2 ), .ZN(
        addr_to_iram[29]) );
  TINV_X1 U4404 ( .I(n7710), .EN(\pipeline/stageF/PC_reg/N1 ), .ZN(
        addr_to_iram[30]) );
  DFF_X1 \pipeline/EXMEM_stage/Forward_sw1_mux_reg  ( .D(
        \pipeline/EXMEM_stage/N76 ), .CK(Clk), .Q(\pipeline/Forward_sw1_mux ), 
        .QN(n17380) );
  DFF_X1 \pipeline/MEMWB_Stage/RegDst_Addr_out_MEMWB_reg[4]  ( .D(
        \pipeline/MEMWB_Stage/N47 ), .CK(Clk), .Q(\pipeline/RegDst_to_WB[4] ), 
        .QN(n17386) );
  DFF_X1 \pipeline/MEMWB_Stage/RegDst_Addr_out_MEMWB_reg[1]  ( .D(
        \pipeline/MEMWB_Stage/N44 ), .CK(Clk), .Q(\pipeline/RegDst_to_WB[1] ), 
        .QN(n17304) );
  DFF_X1 \pipeline/IDEX_Stage/Reg2_Addr_out_IDEX_reg[1]  ( .D(
        \pipeline/IDEX_Stage/N204 ), .CK(Clk), .Q(
        \pipeline/Reg2_Addr_to_exe [1]) );
  DFF_X1 \pipeline/IDEX_Stage/Reg1_Addr_out_IDEX_reg[0]  ( .D(
        \pipeline/IDEX_Stage/N198 ), .CK(Clk), .Q(
        \pipeline/Reg1_Addr_to_exe [0]) );
  DFF_X1 \pipeline/IFID_stage/PC_out_IFID_reg[27]  ( .D(n3909), .CK(Clk), .Q(
        \pipeline/nextPC_IFID_DEC[27] ), .QN(n17469) );
  DFF_X1 \pipeline/IFID_stage/PC_out_IFID_reg[26]  ( .D(n3907), .CK(Clk), .Q(
        \pipeline/nextPC_IFID_DEC[26] ), .QN(n17466) );
  DFF_X1 \pipeline/IFID_stage/PC_out_IFID_reg[25]  ( .D(n3905), .CK(Clk), .Q(
        \pipeline/nextPC_IFID_DEC[25] ), .QN(n17451) );
  DFF_X1 \pipeline/IFID_stage/PC_out_IFID_reg[24]  ( .D(n3903), .CK(Clk), .Q(
        \pipeline/nextPC_IFID_DEC[24] ), .QN(n17465) );
  DFF_X1 \pipeline/IFID_stage/PC_out_IFID_reg[23]  ( .D(n3901), .CK(Clk), .Q(
        \pipeline/nextPC_IFID_DEC[23] ), .QN(n17435) );
  DFF_X1 \pipeline/IFID_stage/PC_out_IFID_reg[22]  ( .D(n3899), .CK(Clk), .Q(
        \pipeline/nextPC_IFID_DEC[22] ), .QN(n17464) );
  DFF_X1 \pipeline/IFID_stage/PC_out_IFID_reg[21]  ( .D(n3897), .CK(Clk), .Q(
        \pipeline/nextPC_IFID_DEC[21] ), .QN(n17448) );
  DFF_X1 \pipeline/IFID_stage/PC_out_IFID_reg[20]  ( .D(n3895), .CK(Clk), .Q(
        \pipeline/nextPC_IFID_DEC[20] ), .QN(n17463) );
  DFF_X1 \pipeline/IFID_stage/PC_out_IFID_reg[19]  ( .D(n3893), .CK(Clk), .Q(
        \pipeline/nextPC_IFID_DEC[19] ), .QN(n17438) );
  DFF_X1 \pipeline/IFID_stage/PC_out_IFID_reg[18]  ( .D(n3891), .CK(Clk), .Q(
        \pipeline/nextPC_IFID_DEC[18] ), .QN(n17462) );
  DFF_X1 \pipeline/IFID_stage/PC_out_IFID_reg[17]  ( .D(n3889), .CK(Clk), .Q(
        \pipeline/nextPC_IFID_DEC[17] ), .QN(n17443) );
  DFF_X1 \pipeline/IFID_stage/PC_out_IFID_reg[15]  ( .D(n3887), .CK(Clk), .Q(
        \pipeline/nextPC_IFID_DEC[15] ), .QN(n17453) );
  DFF_X1 \pipeline/IFID_stage/PC_out_IFID_reg[14]  ( .D(n3885), .CK(Clk), .Q(
        \pipeline/nextPC_IFID_DEC[14] ), .QN(n17460) );
  DFF_X1 \pipeline/IFID_stage/PC_out_IFID_reg[13]  ( .D(n3883), .CK(Clk), .Q(
        \pipeline/nextPC_IFID_DEC[13] ), .QN(n17442) );
  DFF_X1 \pipeline/IFID_stage/PC_out_IFID_reg[12]  ( .D(n3861), .CK(Clk), .Q(
        \pipeline/nextPC_IFID_DEC[12] ), .QN(n17459) );
  DFF_X1 \pipeline/IFID_stage/PC_out_IFID_reg[11]  ( .D(n3867), .CK(Clk), .Q(
        \pipeline/nextPC_IFID_DEC[11] ), .QN(n17441) );
  DFF_X1 \pipeline/IFID_stage/PC_out_IFID_reg[10]  ( .D(n3863), .CK(Clk), .Q(
        \pipeline/nextPC_IFID_DEC[10] ), .QN(n17458) );
  DFF_X1 \pipeline/IFID_stage/PC_out_IFID_reg[9]  ( .D(n3865), .CK(Clk), .Q(
        \pipeline/nextPC_IFID_DEC[9] ), .QN(n17436) );
  DFF_X1 \pipeline/IFID_stage/PC_out_IFID_reg[8]  ( .D(n3881), .CK(Clk), .Q(
        \pipeline/nextPC_IFID_DEC[8] ), .QN(n17457) );
  DFF_X1 \pipeline/IFID_stage/PC_out_IFID_reg[7]  ( .D(n3875), .CK(Clk), .Q(
        \pipeline/nextPC_IFID_DEC[7] ), .QN(n17468) );
  DFF_X1 \pipeline/IFID_stage/PC_out_IFID_reg[6]  ( .D(n3869), .CK(Clk), .Q(
        \pipeline/nextPC_IFID_DEC[6] ), .QN(n17456) );
  DFF_X1 \pipeline/IFID_stage/PC_out_IFID_reg[5]  ( .D(n3871), .CK(Clk), .Q(
        \pipeline/nextPC_IFID_DEC[5] ), .QN(n17454) );
  DFF_X1 \pipeline/IFID_stage/PC_out_IFID_reg[4]  ( .D(n3873), .CK(Clk), .Q(
        \pipeline/nextPC_IFID_DEC[4] ), .QN(n17455) );
  DFF_X1 \pipeline/IFID_stage/PC_out_IFID_reg[3]  ( .D(n3877), .CK(Clk), .Q(
        \pipeline/nextPC_IFID_DEC[3] ), .QN(n17439) );
  DFF_X1 \pipeline/IFID_stage/PC_out_IFID_reg[2]  ( .D(n3859), .CK(Clk), .Q(
        \pipeline/nextPC_IFID_DEC[2] ), .QN(n17470) );
  DFF_X1 \pipeline/IFID_stage/Instr_out_IFID_reg[31]  ( .D(n3957), .CK(Clk), 
        .Q(\pipeline/inst_IFID_DEC[31] ), .QN(n17532) );
  DFF_X1 \pipeline/IFID_stage/Instr_out_IFID_reg[23]  ( .D(n3965), .CK(Clk), 
        .Q(\pipeline/stageD/offset_jump_sign_ext [23]), .QN(n17383) );
  DFF_X1 \pipeline/EXMEM_stage/ALUres_MEMaddr_out_EXMEM_reg[11]  ( .D(
        \pipeline/EXMEM_stage/N18 ), .CK(Clk), .Q(
        \pipeline/Alu_Out_Addr_to_mem[11] ) );
  DFF_X1 \pipeline/EXMEM_stage/ALUres_MEMaddr_out_EXMEM_reg[9]  ( .D(
        \pipeline/EXMEM_stage/N16 ), .CK(Clk), .Q(
        \pipeline/Alu_Out_Addr_to_mem[9] ) );
  DFF_X1 \pipeline/EXMEM_stage/ALUres_MEMaddr_out_EXMEM_reg[10]  ( .D(
        \pipeline/EXMEM_stage/N17 ), .CK(Clk), .Q(
        \pipeline/Alu_Out_Addr_to_mem[10] ) );
  DFF_X1 \pipeline/EXMEM_stage/ALUres_MEMaddr_out_EXMEM_reg[8]  ( .D(
        \pipeline/EXMEM_stage/N15 ), .CK(Clk), .Q(
        \pipeline/Alu_Out_Addr_to_mem[8] ) );
  DFF_X1 \pipeline/EXMEM_stage/ALUres_MEMaddr_out_EXMEM_reg[2]  ( .D(
        \pipeline/EXMEM_stage/N9 ), .CK(Clk), .Q(
        \pipeline/Alu_Out_Addr_to_mem[2] ), .QN(n17398) );
  DFF_X1 \pipeline/IFID_stage/PC_out_IFID_reg[28]  ( .D(n3911), .CK(Clk), .Q(
        \pipeline/nextPC_IFID_DEC[28] ), .QN(n17467) );
  DFF_X1 \pipeline/EXMEM_stage/ALUres_MEMaddr_out_EXMEM_reg[1]  ( .D(
        \pipeline/EXMEM_stage/N8 ), .CK(Clk), .Q(
        \pipeline/Alu_Out_Addr_to_mem[1] ), .QN(n17397) );
  DFF_X1 \pipeline/EXMEM_stage/ALUres_MEMaddr_out_EXMEM_reg[5]  ( .D(
        \pipeline/EXMEM_stage/N12 ), .CK(Clk), .Q(
        \pipeline/Alu_Out_Addr_to_mem[5] ) );
  DFF_X1 \pipeline/EXMEM_stage/ALUres_MEMaddr_out_EXMEM_reg[6]  ( .D(
        \pipeline/EXMEM_stage/N13 ), .CK(Clk), .Q(
        \pipeline/Alu_Out_Addr_to_mem[6] ) );
  DFF_X1 \pipeline/EXMEM_stage/ALUres_MEMaddr_out_EXMEM_reg[4]  ( .D(
        \pipeline/EXMEM_stage/N11 ), .CK(Clk), .Q(
        \pipeline/Alu_Out_Addr_to_mem[4] ) );
  DFF_X1 \pipeline/EXMEM_stage/ALUres_MEMaddr_out_EXMEM_reg[3]  ( .D(
        \pipeline/EXMEM_stage/N10 ), .CK(Clk), .Q(
        \pipeline/Alu_Out_Addr_to_mem[3] ) );
  DFF_X1 \pipeline/EXMEM_stage/ALUres_MEMaddr_out_EXMEM_reg[13]  ( .D(
        \pipeline/EXMEM_stage/N20 ), .CK(Clk), .Q(
        \pipeline/Alu_Out_Addr_to_mem[13] ) );
  DFF_X1 \pipeline/IFID_stage/PC_out_IFID_reg[29]  ( .D(n3856), .CK(Clk), .Q(
        \pipeline/nextPC_IFID_DEC[29] ), .QN(n17452) );
  DFF_X1 \pipeline/EXMEM_stage/ALUres_MEMaddr_out_EXMEM_reg[14]  ( .D(
        \pipeline/EXMEM_stage/N21 ), .CK(Clk), .Q(
        \pipeline/Alu_Out_Addr_to_mem[14] ) );
  DFF_X1 \pipeline/IFID_stage/PC_out_IFID_reg[30]  ( .D(n3855), .CK(Clk), .Q(
        \pipeline/nextPC_IFID_DEC[30] ), .QN(n17471) );
  DFF_X1 \pipeline/EXMEM_stage/ALUres_MEMaddr_out_EXMEM_reg[16]  ( .D(
        \pipeline/EXMEM_stage/N23 ), .CK(Clk), .Q(
        \pipeline/Alu_Out_Addr_to_mem[16] ) );
  DFF_X1 \pipeline/EXMEM_stage/ALUres_MEMaddr_out_EXMEM_reg[15]  ( .D(
        \pipeline/EXMEM_stage/N22 ), .CK(Clk), .Q(
        \pipeline/Alu_Out_Addr_to_mem[15] ) );
  DFF_X1 \pipeline/EXMEM_stage/ALUres_MEMaddr_out_EXMEM_reg[17]  ( .D(
        \pipeline/EXMEM_stage/N24 ), .CK(Clk), .Q(
        \pipeline/Alu_Out_Addr_to_mem[17] ) );
  DFF_X1 \pipeline/EXMEM_stage/ALUres_MEMaddr_out_EXMEM_reg[22]  ( .D(
        \pipeline/EXMEM_stage/N29 ), .CK(Clk), .Q(
        \pipeline/Alu_Out_Addr_to_mem[22] ) );
  DFF_X1 \pipeline/EXMEM_stage/ALUres_MEMaddr_out_EXMEM_reg[20]  ( .D(
        \pipeline/EXMEM_stage/N27 ), .CK(Clk), .Q(
        \pipeline/Alu_Out_Addr_to_mem[20] ) );
  DFF_X1 \pipeline/EXMEM_stage/ALUres_MEMaddr_out_EXMEM_reg[21]  ( .D(
        \pipeline/EXMEM_stage/N28 ), .CK(Clk), .Q(
        \pipeline/Alu_Out_Addr_to_mem[21] ) );
  DFF_X1 \pipeline/EXMEM_stage/ALUres_MEMaddr_out_EXMEM_reg[19]  ( .D(
        \pipeline/EXMEM_stage/N26 ), .CK(Clk), .Q(
        \pipeline/Alu_Out_Addr_to_mem[19] ) );
  DFF_X1 \pipeline/EXMEM_stage/ALUres_MEMaddr_out_EXMEM_reg[23]  ( .D(
        \pipeline/EXMEM_stage/N30 ), .CK(Clk), .Q(
        \pipeline/Alu_Out_Addr_to_mem[23] ) );
  DFF_X1 \pipeline/EXMEM_stage/ALUres_MEMaddr_out_EXMEM_reg[18]  ( .D(
        \pipeline/EXMEM_stage/N25 ), .CK(Clk), .Q(
        \pipeline/Alu_Out_Addr_to_mem[18] ) );
  DFF_X1 \pipeline/EXMEM_stage/ALUres_MEMaddr_out_EXMEM_reg[25]  ( .D(
        \pipeline/EXMEM_stage/N32 ), .CK(Clk), .Q(
        \pipeline/Alu_Out_Addr_to_mem[25] ) );
  DFF_X1 \pipeline/EXMEM_stage/ALUres_MEMaddr_out_EXMEM_reg[26]  ( .D(
        \pipeline/EXMEM_stage/N33 ), .CK(Clk), .Q(
        \pipeline/Alu_Out_Addr_to_mem[26] ) );
  DFF_X1 \pipeline/EXMEM_stage/ALUres_MEMaddr_out_EXMEM_reg[24]  ( .D(
        \pipeline/EXMEM_stage/N31 ), .CK(Clk), .Q(
        \pipeline/Alu_Out_Addr_to_mem[24] ) );
  DFF_X1 \pipeline/EXMEM_stage/ALUres_MEMaddr_out_EXMEM_reg[27]  ( .D(
        \pipeline/EXMEM_stage/N34 ), .CK(Clk), .Q(
        \pipeline/Alu_Out_Addr_to_mem[27] ) );
  DFF_X1 \pipeline/EXMEM_stage/ALUres_MEMaddr_out_EXMEM_reg[28]  ( .D(
        \pipeline/EXMEM_stage/N35 ), .CK(Clk), .Q(
        \pipeline/Alu_Out_Addr_to_mem[28] ) );
  DFF_X1 \pipeline/EXMEM_stage/ALUres_MEMaddr_out_EXMEM_reg[29]  ( .D(
        \pipeline/EXMEM_stage/N36 ), .CK(Clk), .Q(
        \pipeline/Alu_Out_Addr_to_mem[29] ) );
  DFF_X1 \pipeline/EXMEM_stage/ALUres_MEMaddr_out_EXMEM_reg[30]  ( .D(
        \pipeline/EXMEM_stage/N37 ), .CK(Clk), .Q(
        \pipeline/Alu_Out_Addr_to_mem[30] ) );
  DFF_X1 \pipeline/EXMEM_stage/ALUres_MEMaddr_out_EXMEM_reg[31]  ( .D(
        \pipeline/EXMEM_stage/N38 ), .CK(Clk), .Q(
        \pipeline/Alu_Out_Addr_to_mem[31] ) );
  DFF_X1 \pipeline/IFID_stage/PC_out_IFID_reg[1]  ( .D(n3857), .CK(Clk), .Q(
        \pipeline/nextPC_IFID_DEC[1] ), .QN(n17446) );
  DFF_X1 \pipeline/IDEX_Stage/Reg2_Addr_out_IDEX_reg[4]  ( .D(
        \pipeline/IDEX_Stage/N207 ), .CK(Clk), .Q(
        \pipeline/Reg2_Addr_to_exe [4]) );
  DFF_X1 \pipeline/EXMEM_stage/RegDst_Addr_out_EXMEM_reg[0]  ( .D(
        \pipeline/EXMEM_stage/N71 ), .CK(Clk), .Q(\pipeline/regDst_to_mem[0] ), 
        .QN(n17644) );
  DFF_X1 \pipeline/EXMEM_stage/RegDst_Addr_out_EXMEM_reg[3]  ( .D(
        \pipeline/EXMEM_stage/N74 ), .CK(Clk), .Q(\pipeline/regDst_to_mem[3] ), 
        .QN(n17340) );
  DFF_X1 \pipeline/EXMEM_stage/RegDst_Addr_out_EXMEM_reg[4]  ( .D(
        \pipeline/EXMEM_stage/N75 ), .CK(Clk), .Q(\pipeline/regDst_to_mem[4] ), 
        .QN(n17393) );
  DFF_X1 \pipeline/EXMEM_stage/ALUres_MEMaddr_out_EXMEM_reg[0]  ( .D(
        \pipeline/EXMEM_stage/N7 ), .CK(Clk), .Q(
        \pipeline/Alu_Out_Addr_to_mem[0] ) );
  DFF_X1 \pipeline/IFID_stage/Instr_out_IFID_reg[4]  ( .D(n3983), .CK(Clk), 
        .Q(\pipeline/stageD/offset_to_jump_temp [4]), .QN(n17412) );
  NAND3_X1 U11979 ( .A1(n13980), .A2(n17704), .A3(n13984), .ZN(
        \pipeline/cu_pipeline/N107 ) );
  NAND3_X1 U11980 ( .A1(n14028), .A2(n14019), .A3(n14029), .ZN(n14027) );
  NAND3_X1 U11981 ( .A1(\pipeline/inst_IFID_DEC[29] ), .A2(n13995), .A3(n17348), .ZN(n14035) );
  NAND3_X1 U11982 ( .A1(n14005), .A2(n14044), .A3(n14032), .ZN(n14021) );
  NAND3_X1 U11983 ( .A1(n14049), .A2(n14000), .A3(n17382), .ZN(n14048) );
  NAND3_X1 U11984 ( .A1(n14000), .A2(n17348), .A3(\pipeline/inst_IFID_DEC[29] ), .ZN(n14070) );
  NAND3_X1 U11985 ( .A1(\pipeline/WB_controls_in_MEMWB[1] ), .A2(
        \pipeline/MEM_controls_in_MEM[1] ), .A3(n14090), .ZN(n14089) );
  NAND3_X1 U11986 ( .A1(\pipeline/WB_controls_in_EXMEM[1] ), .A2(
        \pipeline/MEM_controls_in_EXMEM[1] ), .A3(n14095), .ZN(n14086) );
  XOR2_X1 U11987 ( .A(n17384), .B(n14100), .Z(n14099) );
  XOR2_X1 U11988 ( .A(n17328), .B(n14101), .Z(n14097) );
  XOR2_X1 U11993 ( .A(n17383), .B(n14113), .Z(n14098) );
  NAND3_X1 U11994 ( .A1(\pipeline/WB_controls_in_EXMEM[1] ), .A2(
        \pipeline/MEM_controls_in_EXMEM[1] ), .A3(n13983), .ZN(n14094) );
  NAND3_X1 U11995 ( .A1(\pipeline/cu_pipeline/N89 ), .A2(n17428), .A3(n17361), 
        .ZN(n14174) );
  NAND3_X1 U11996 ( .A1(\pipeline/stageD/offset_to_jump_temp [5]), .A2(n14067), 
        .A3(n17406), .ZN(n14066) );
  NAND3_X1 U11997 ( .A1(\pipeline/inst_IFID_DEC[29] ), .A2(n14049), .A3(n17313), .ZN(n14058) );
  NAND3_X1 U11998 ( .A1(\pipeline/inst_IFID_DEC[27] ), .A2(n14001), .A3(n17347), .ZN(n14029) );
  NAND3_X1 U11999 ( .A1(\pipeline/inst_IFID_DEC[31] ), .A2(n14084), .A3(n17348), .ZN(n14169) );
  NAND3_X1 U12000 ( .A1(n14241), .A2(n14242), .A3(n14243), .ZN(n14201) );
  NAND3_X1 U12001 ( .A1(n14268), .A2(n14269), .A3(n14270), .ZN(n14252) );
  NAND3_X1 U12002 ( .A1(n14288), .A2(n14289), .A3(n14290), .ZN(n14272) );
  NAND3_X1 U12003 ( .A1(n14308), .A2(n14309), .A3(n14310), .ZN(n14292) );
  NAND3_X1 U12004 ( .A1(n14328), .A2(n14329), .A3(n14330), .ZN(n14312) );
  NAND3_X1 U12005 ( .A1(n14348), .A2(n14349), .A3(n14350), .ZN(n14332) );
  NAND3_X1 U12006 ( .A1(n14368), .A2(n14369), .A3(n14370), .ZN(n14352) );
  NAND3_X1 U12007 ( .A1(n14388), .A2(n14389), .A3(n14390), .ZN(n14372) );
  NAND3_X1 U12008 ( .A1(n14408), .A2(n14409), .A3(n14410), .ZN(n14392) );
  NAND3_X1 U12009 ( .A1(n14428), .A2(n14429), .A3(n14430), .ZN(n14412) );
  NAND3_X1 U12010 ( .A1(n14448), .A2(n14449), .A3(n14450), .ZN(n14432) );
  NAND3_X1 U12011 ( .A1(n14468), .A2(n14469), .A3(n14470), .ZN(n14452) );
  NAND3_X1 U12012 ( .A1(n14488), .A2(n14489), .A3(n14490), .ZN(n14472) );
  NAND3_X1 U12013 ( .A1(n14508), .A2(n14509), .A3(n14510), .ZN(n14492) );
  NAND3_X1 U12014 ( .A1(n14528), .A2(n14529), .A3(n14530), .ZN(n14512) );
  NAND3_X1 U12015 ( .A1(n14548), .A2(n14549), .A3(n14550), .ZN(n14532) );
  NAND3_X1 U12016 ( .A1(n14568), .A2(n14569), .A3(n14570), .ZN(n14552) );
  NAND3_X1 U12017 ( .A1(n14588), .A2(n14589), .A3(n14590), .ZN(n14572) );
  NAND3_X1 U12018 ( .A1(n14608), .A2(n14609), .A3(n14610), .ZN(n14592) );
  NAND3_X1 U12019 ( .A1(n14628), .A2(n14629), .A3(n14630), .ZN(n14612) );
  NAND3_X1 U12020 ( .A1(n14648), .A2(n14649), .A3(n14650), .ZN(n14632) );
  NAND3_X1 U12021 ( .A1(n14668), .A2(n14669), .A3(n14670), .ZN(n14652) );
  NAND3_X1 U12022 ( .A1(n14688), .A2(n14689), .A3(n14690), .ZN(n14672) );
  NAND3_X1 U12023 ( .A1(n14708), .A2(n14709), .A3(n14710), .ZN(n14692) );
  NAND3_X1 U12024 ( .A1(n14728), .A2(n14729), .A3(n14730), .ZN(n14712) );
  NAND3_X1 U12025 ( .A1(n14748), .A2(n14749), .A3(n14750), .ZN(n14732) );
  NAND3_X1 U12026 ( .A1(n14768), .A2(n14769), .A3(n14770), .ZN(n14752) );
  NAND3_X1 U12027 ( .A1(n14788), .A2(n14789), .A3(n14790), .ZN(n14772) );
  NAND3_X1 U12028 ( .A1(n14808), .A2(n14809), .A3(n14810), .ZN(n14792) );
  NAND3_X1 U12029 ( .A1(n14828), .A2(n14829), .A3(n14830), .ZN(n14812) );
  NAND3_X1 U12030 ( .A1(n14848), .A2(n14849), .A3(n14850), .ZN(n14832) );
  NAND3_X1 U12031 ( .A1(\pipeline/stageD/offset_jump_sign_ext [16]), .A2(
        n17407), .A3(n17349), .ZN(n14861) );
  NAND3_X1 U12032 ( .A1(\pipeline/stageD/offset_jump_sign_ext [19]), .A2(
        \pipeline/stageD/offset_jump_sign_ext [16]), .A3(n17407), .ZN(n14867)
         );
  NAND3_X1 U12033 ( .A1(\pipeline/stageD/offset_jump_sign_ext [19]), .A2(
        n17407), .A3(n17316), .ZN(n14866) );
  NAND3_X1 U12034 ( .A1(\pipeline/stageD/offset_jump_sign_ext [20]), .A2(
        n17349), .A3(n17316), .ZN(n14872) );
  NAND3_X1 U12035 ( .A1(\pipeline/stageD/offset_jump_sign_ext [20]), .A2(
        \pipeline/stageD/offset_jump_sign_ext [16]), .A3(n17349), .ZN(n14873)
         );
  NAND3_X1 U12036 ( .A1(n14880), .A2(n14881), .A3(n14882), .ZN(n14852) );
  NAND3_X1 U12037 ( .A1(n17407), .A2(n17349), .A3(n17316), .ZN(n14862) );
  NAND3_X1 U12038 ( .A1(\pipeline/stageD/offset_jump_sign_ext [19]), .A2(
        \pipeline/stageD/offset_jump_sign_ext [20]), .A3(n17316), .ZN(n14878)
         );
  NAND3_X1 U12039 ( .A1(\pipeline/stageD/offset_jump_sign_ext [20]), .A2(
        \pipeline/stageD/offset_jump_sign_ext [19]), .A3(
        \pipeline/stageD/offset_jump_sign_ext [16]), .ZN(n14879) );
  NAND3_X1 U12040 ( .A1(n14952), .A2(n12649), .A3(n17740), .ZN(n14951) );
  NAND3_X1 U12041 ( .A1(n14958), .A2(n14959), .A3(n14960), .ZN(n14957) );
  OAI33_X1 U12042 ( .A1(n17074), .A2(n14967), .A3(n12649), .B1(n17740), .B2(
        n14968), .B3(n17091), .ZN(n14956) );
  NAND3_X1 U12043 ( .A1(n17103), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[1] ), .A3(n14954), .ZN(
        n14972) );
  NAND3_X1 U12044 ( .A1(n14977), .A2(n14978), .A3(n14979), .ZN(n14976) );
  MUX2_X1 U12045 ( .A(n13934), .B(n13929), .S(n17430), .Z(n14120) );
  NAND3_X1 U12046 ( .A1(n17104), .A2(n15133), .A3(n14954), .ZN(n15131) );
  OAI33_X1 U12047 ( .A1(n15133), .A2(n17679), .A3(
        \pipeline/stageE/EXE_ALU/alu_shift/N136 ), .B1(n15134), .B2(n14968), 
        .B3(n17104), .ZN(n15126) );
  NAND3_X1 U12050 ( .A1(\pipeline/stageE/EXE_ALU/alu_shift/N136 ), .A2(n14952), 
        .A3(n15134), .ZN(n15124) );
  NAND3_X1 U12051 ( .A1(n14952), .A2(\pipeline/stageE/input1_to_ALU [30]), 
        .A3(n15150), .ZN(n15149) );
  NAND3_X1 U12052 ( .A1(n15154), .A2(n15155), .A3(n15156), .ZN(n15153) );
  OAI33_X1 U12053 ( .A1(n15157), .A2(n17678), .A3(
        \pipeline/stageE/input1_to_ALU [30]), .B1(n15150), .B2(n14968), .B3(
        n17083), .ZN(n15152) );
  XOR2_X1 U12054 ( .A(n15159), .B(n15160), .Z(n15009) );
  NAND3_X1 U12055 ( .A1(n14952), .A2(\pipeline/stageE/input1_to_ALU [29]), 
        .A3(n15169), .ZN(n15168) );
  NAND3_X1 U12056 ( .A1(n15173), .A2(n15174), .A3(n15175), .ZN(n15172) );
  OAI33_X1 U12057 ( .A1(n15176), .A2(n14967), .A3(
        \pipeline/stageE/input1_to_ALU [29]), .B1(n15169), .B2(n14968), .B3(
        n17094), .ZN(n15171) );
  NAND3_X1 U12058 ( .A1(n14952), .A2(\pipeline/stageE/input1_to_ALU [28]), 
        .A3(n15182), .ZN(n15181) );
  NAND3_X1 U12059 ( .A1(n15186), .A2(n15187), .A3(n15188), .ZN(n15185) );
  OAI33_X1 U12060 ( .A1(n15189), .A2(n17679), .A3(
        \pipeline/stageE/input1_to_ALU [28]), .B1(n15182), .B2(n14968), .B3(
        n17093), .ZN(n15184) );
  NAND3_X1 U12061 ( .A1(n17078), .A2(n15201), .A3(n14954), .ZN(n15199) );
  OAI33_X1 U12062 ( .A1(n15201), .A2(n17678), .A3(
        \pipeline/stageE/input1_to_ALU [27]), .B1(n15202), .B2(n14968), .B3(
        n17078), .ZN(n15194) );
  NAND3_X1 U12064 ( .A1(\pipeline/stageE/input1_to_ALU [27]), .A2(n14952), 
        .A3(n15202), .ZN(n15192) );
  NAND3_X1 U12065 ( .A1(n17086), .A2(n15215), .A3(n14954), .ZN(n15213) );
  OAI33_X1 U12066 ( .A1(n15215), .A2(n14967), .A3(
        \pipeline/stageE/input1_to_ALU [26]), .B1(n15216), .B2(n14968), .B3(
        n17086), .ZN(n15208) );
  NAND3_X1 U12067 ( .A1(\pipeline/stageE/input1_to_ALU [26]), .A2(n14952), 
        .A3(n15216), .ZN(n15206) );
  NAND3_X1 U12068 ( .A1(n14952), .A2(n17159), .A3(n15224), .ZN(n15223) );
  NAND3_X1 U12069 ( .A1(n15228), .A2(n15229), .A3(n15230), .ZN(n15227) );
  OAI33_X1 U12070 ( .A1(n15231), .A2(n17679), .A3(n17159), .B1(n15224), .B2(
        n14968), .B3(n17115), .ZN(n15226) );
  NAND3_X1 U12071 ( .A1(n17117), .A2(n15245), .A3(n14954), .ZN(n15243) );
  OAI33_X1 U12072 ( .A1(n15245), .A2(n17678), .A3(n17158), .B1(n15246), .B2(
        n14968), .B3(n17117), .ZN(n15238) );
  XOR2_X1 U12073 ( .A(n15247), .B(n15248), .Z(n15013) );
  NAND3_X1 U12074 ( .A1(n17158), .A2(n14952), .A3(n15246), .ZN(n15236) );
  NAND3_X1 U12075 ( .A1(n17092), .A2(n15260), .A3(n17677), .ZN(n15258) );
  OAI33_X1 U12076 ( .A1(n15260), .A2(n14967), .A3(
        \pipeline/stageE/input1_to_ALU [23]), .B1(n15261), .B2(n14968), .B3(
        n17092), .ZN(n15253) );
  XOR2_X1 U12077 ( .A(n15262), .B(n15263), .Z(n15022) );
  NAND3_X1 U12078 ( .A1(\pipeline/stageE/input1_to_ALU [23]), .A2(n14952), 
        .A3(n15261), .ZN(n15251) );
  NAND3_X1 U12079 ( .A1(n17116), .A2(n15278), .A3(n17677), .ZN(n15276) );
  OAI33_X1 U12080 ( .A1(n15278), .A2(n17679), .A3(
        \pipeline/stageE/input1_to_ALU [22]), .B1(n15279), .B2(n14968), .B3(
        n17116), .ZN(n15271) );
  NAND3_X1 U12081 ( .A1(\pipeline/stageE/input1_to_ALU [22]), .A2(n14952), 
        .A3(n15279), .ZN(n15269) );
  NAND3_X1 U12082 ( .A1(n14952), .A2(\pipeline/stageE/input1_to_ALU [21]), 
        .A3(n15285), .ZN(n15284) );
  NAND3_X1 U12083 ( .A1(n15289), .A2(n15290), .A3(n15291), .ZN(n15288) );
  OAI33_X1 U12084 ( .A1(n15292), .A2(n17678), .A3(
        \pipeline/stageE/input1_to_ALU [21]), .B1(n15285), .B2(n14968), .B3(
        n17084), .ZN(n15287) );
  XOR2_X1 U12085 ( .A(n15294), .B(n15295), .Z(n15017) );
  NAND3_X1 U12086 ( .A1(n17118), .A2(n15311), .A3(n17677), .ZN(n15309) );
  OAI33_X1 U12087 ( .A1(n15311), .A2(n14967), .A3(n17157), .B1(n15312), .B2(
        n14968), .B3(n17118), .ZN(n15304) );
  NAND3_X1 U12088 ( .A1(n17157), .A2(n14952), .A3(n15312), .ZN(n15302) );
  NAND3_X1 U12089 ( .A1(n17097), .A2(n15330), .A3(n17677), .ZN(n15328) );
  OAI33_X1 U12090 ( .A1(n15330), .A2(n17679), .A3(
        \pipeline/stageE/input1_to_ALU [19]), .B1(n15331), .B2(n14968), .B3(
        n17097), .ZN(n15323) );
  XOR2_X1 U12091 ( .A(n15332), .B(n15333), .Z(n15023) );
  XOR2_X1 U12092 ( .A(n15334), .B(n17097), .Z(n15333) );
  NAND3_X1 U12093 ( .A1(\pipeline/stageE/input1_to_ALU [19]), .A2(n14952), 
        .A3(n15331), .ZN(n15321) );
  NAND3_X1 U12094 ( .A1(n17096), .A2(n15345), .A3(n17677), .ZN(n15343) );
  OAI33_X1 U12095 ( .A1(n15345), .A2(n17678), .A3(
        \pipeline/stageE/input1_to_ALU [18]), .B1(n15346), .B2(n14968), .B3(
        n17096), .ZN(n15338) );
  NAND3_X1 U12097 ( .A1(\pipeline/stageE/input1_to_ALU [18]), .A2(n14952), 
        .A3(n15346), .ZN(n15336) );
  NAND3_X1 U12098 ( .A1(n17079), .A2(n15362), .A3(n17677), .ZN(n15360) );
  OAI33_X1 U12099 ( .A1(n15362), .A2(n14967), .A3(
        \pipeline/stageE/input1_to_ALU [17]), .B1(n15363), .B2(n14968), .B3(
        n17079), .ZN(n15355) );
  NAND3_X1 U12101 ( .A1(\pipeline/stageE/input1_to_ALU [17]), .A2(n14952), 
        .A3(n15363), .ZN(n15353) );
  NAND3_X1 U12102 ( .A1(n14952), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/A[16] ), .A3(n15372), .ZN(
        n15371) );
  NAND3_X1 U12103 ( .A1(n15376), .A2(n15377), .A3(n15378), .ZN(n15375) );
  OAI33_X1 U12104 ( .A1(n15379), .A2(n17679), .A3(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/A[16] ), .B1(n15372), .B2(
        n14968), .B3(n17738), .ZN(n15374) );
  XOR2_X1 U12105 ( .A(n15381), .B(n15368), .Z(n15032) );
  NAND3_X1 U12106 ( .A1(n14952), .A2(\pipeline/stageE/input1_to_ALU [15]), 
        .A3(n15386), .ZN(n15385) );
  NAND3_X1 U12107 ( .A1(n15390), .A2(n15391), .A3(n15392), .ZN(n15389) );
  OAI33_X1 U12108 ( .A1(n15393), .A2(n17678), .A3(
        \pipeline/stageE/input1_to_ALU [15]), .B1(n15386), .B2(n14968), .B3(
        n17101), .ZN(n15388) );
  XOR2_X1 U12109 ( .A(n15395), .B(n15396), .Z(n15029) );
  XOR2_X1 U12110 ( .A(n17101), .B(n15397), .Z(n15396) );
  NAND3_X1 U12111 ( .A1(n17100), .A2(n15410), .A3(n17677), .ZN(n15408) );
  OAI33_X1 U12112 ( .A1(n15410), .A2(n14967), .A3(
        \pipeline/stageE/input1_to_ALU [14]), .B1(n15411), .B2(n14968), .B3(
        n17100), .ZN(n15403) );
  XOR2_X1 U12113 ( .A(n15399), .B(n15412), .Z(n15027) );
  NAND3_X1 U12114 ( .A1(\pipeline/stageE/input1_to_ALU [14]), .A2(n14952), 
        .A3(n15411), .ZN(n15401) );
  NAND3_X1 U12115 ( .A1(n15425), .A2(n15426), .A3(n17677), .ZN(n15424) );
  OAI33_X1 U12116 ( .A1(n15426), .A2(n17679), .A3(n17160), .B1(n15427), .B2(
        n14968), .B3(n15425), .ZN(n15419) );
  XOR2_X1 U12117 ( .A(n15428), .B(n15415), .Z(n15033) );
  NAND3_X1 U12118 ( .A1(n17160), .A2(n14952), .A3(n15427), .ZN(n15417) );
  NAND3_X1 U12119 ( .A1(n14952), .A2(\pipeline/stageE/input1_to_ALU [12]), 
        .A3(n15435), .ZN(n15434) );
  NAND3_X1 U12120 ( .A1(n15439), .A2(n15440), .A3(n15441), .ZN(n15438) );
  OAI33_X1 U12121 ( .A1(n15442), .A2(n17678), .A3(
        \pipeline/stageE/input1_to_ALU [12]), .B1(n15435), .B2(n14968), .B3(
        n17080), .ZN(n15437) );
  XOR2_X1 U12122 ( .A(n15444), .B(n15429), .Z(n15030) );
  NAND3_X1 U12123 ( .A1(n14952), .A2(\pipeline/stageE/input1_to_ALU [11]), 
        .A3(n15449), .ZN(n15448) );
  NAND3_X1 U12124 ( .A1(n15453), .A2(n15454), .A3(n15455), .ZN(n15452) );
  OAI33_X1 U12125 ( .A1(n15456), .A2(n14967), .A3(
        \pipeline/stageE/input1_to_ALU [11]), .B1(n15449), .B2(n14968), .B3(
        n17082), .ZN(n15451) );
  NAND3_X1 U12126 ( .A1(n17085), .A2(n15473), .A3(n14954), .ZN(n15471) );
  OAI33_X1 U12127 ( .A1(n15473), .A2(n17679), .A3(
        \pipeline/stageE/input1_to_ALU [10]), .B1(n15474), .B2(n14968), .B3(
        n17085), .ZN(n15466) );
  XOR2_X1 U12128 ( .A(n15475), .B(n15462), .Z(n15034) );
  NAND3_X1 U12129 ( .A1(\pipeline/stageE/input1_to_ALU [10]), .A2(n14952), 
        .A3(n15474), .ZN(n15464) );
  NAND3_X1 U12130 ( .A1(n17090), .A2(n15491), .A3(n14954), .ZN(n15489) );
  OAI33_X1 U12131 ( .A1(n15491), .A2(n17678), .A3(
        \pipeline/stageE/input1_to_ALU [9]), .B1(n15492), .B2(n14968), .B3(
        n17090), .ZN(n15484) );
  NAND3_X1 U12132 ( .A1(\pipeline/stageE/input1_to_ALU [9]), .A2(n14952), .A3(
        n15492), .ZN(n15482) );
  NAND3_X1 U12133 ( .A1(n14952), .A2(\pipeline/stageE/input1_to_ALU [8]), .A3(
        n15498), .ZN(n15497) );
  NAND3_X1 U12134 ( .A1(n15502), .A2(n15503), .A3(n15504), .ZN(n15501) );
  OAI33_X1 U12135 ( .A1(n15505), .A2(n14967), .A3(
        \pipeline/stageE/input1_to_ALU [8]), .B1(n15498), .B2(n14968), .B3(
        n17095), .ZN(n15500) );
  XOR2_X1 U12136 ( .A(n15507), .B(n15508), .Z(n15039) );
  NAND3_X1 U12137 ( .A1(n14952), .A2(\pipeline/stageE/input1_to_ALU [7]), .A3(
        n15512), .ZN(n15511) );
  NAND3_X1 U12138 ( .A1(n15516), .A2(n15517), .A3(n15518), .ZN(n15515) );
  OAI33_X1 U12139 ( .A1(n15519), .A2(n17679), .A3(
        \pipeline/stageE/input1_to_ALU [7]), .B1(n15512), .B2(n14968), .B3(
        n17089), .ZN(n15514) );
  NAND3_X1 U12140 ( .A1(n17088), .A2(n15537), .A3(n14954), .ZN(n15535) );
  OAI33_X1 U12141 ( .A1(n15537), .A2(n17678), .A3(
        \pipeline/stageE/input1_to_ALU [6]), .B1(n15538), .B2(n14968), .B3(
        n17088), .ZN(n15530) );
  NAND3_X1 U12142 ( .A1(\pipeline/stageE/input1_to_ALU [6]), .A2(n14952), .A3(
        n15538), .ZN(n15528) );
  NAND3_X1 U12143 ( .A1(n17087), .A2(n15552), .A3(n14954), .ZN(n15550) );
  OAI33_X1 U12144 ( .A1(n15552), .A2(n14967), .A3(
        \pipeline/stageE/input1_to_ALU [5]), .B1(n15553), .B2(n14968), .B3(
        n17087), .ZN(n15545) );
  NAND3_X1 U12145 ( .A1(\pipeline/stageE/input1_to_ALU [5]), .A2(n14952), .A3(
        n15553), .ZN(n15543) );
  NAND3_X1 U12146 ( .A1(n15564), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .A3(n14954), .ZN(
        n15563) );
  OAI33_X1 U12147 ( .A1(\pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .A2(
        n17679), .A3(\pipeline/stageE/input1_to_ALU [4]), .B1(n17737), .B2(
        n14968), .B3(n15564), .ZN(n15558) );
  XOR2_X1 U12148 ( .A(n15566), .B(n15567), .Z(n15041) );
  NAND3_X1 U12149 ( .A1(n14952), .A2(n17739), .A3(
        \pipeline/stageE/input1_to_ALU [3]), .ZN(n15571) );
  NAND3_X1 U12150 ( .A1(n15577), .A2(n15578), .A3(n15579), .ZN(n15576) );
  NAND3_X1 U12151 ( .A1(\pipeline/EXE_controls_in_EXEcute [5]), .A2(
        \pipeline/EXE_controls_in_EXEcute [6]), .A3(n17705), .ZN(n15586) );
  OAI33_X1 U12152 ( .A1(n17077), .A2(n14968), .A3(n17739), .B1(
        \pipeline/stageE/input1_to_ALU [3]), .B2(n17678), .B3(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[3] ), .ZN(n15575) );
  XOR2_X1 U12154 ( .A(n15590), .B(n15591), .Z(n15045) );
  MUX2_X1 U12155 ( .A(n15592), .B(n15593), .S(n17381), .Z(n15591) );
  NAND3_X1 U12156 ( .A1(n15596), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N202 ), 
        .A3(n15050), .ZN(n15595) );
  XOR2_X1 U12157 ( .A(n15598), .B(n17077), .Z(n15590) );
  NAND3_X1 U12158 ( .A1(n15602), .A2(n15603), .A3(n15604), .ZN(n3991) );
  NAND3_X1 U12161 ( .A1(n15689), .A2(n15690), .A3(n15691), .ZN(n3912) );
  NAND3_X1 U12162 ( .A1(n15694), .A2(n15695), .A3(n15696), .ZN(n3910) );
  NAND3_X1 U12163 ( .A1(n15699), .A2(n15700), .A3(n15701), .ZN(n3908) );
  NAND3_X1 U12164 ( .A1(n15704), .A2(n15705), .A3(n15706), .ZN(n3906) );
  NAND3_X1 U12165 ( .A1(n15709), .A2(n15710), .A3(n15711), .ZN(n3904) );
  NAND3_X1 U12166 ( .A1(n15714), .A2(n15715), .A3(n15716), .ZN(n3902) );
  NAND3_X1 U12167 ( .A1(n15719), .A2(n15720), .A3(n15721), .ZN(n3900) );
  NAND3_X1 U12168 ( .A1(n15724), .A2(n15725), .A3(n15726), .ZN(n3898) );
  NAND3_X1 U12169 ( .A1(n15729), .A2(n15730), .A3(n15731), .ZN(n3896) );
  NAND3_X1 U12170 ( .A1(n15734), .A2(n15735), .A3(n15736), .ZN(n3894) );
  NAND3_X1 U12171 ( .A1(n15739), .A2(n15740), .A3(n15741), .ZN(n3892) );
  NAND3_X1 U12172 ( .A1(n15744), .A2(n15745), .A3(n15746), .ZN(n3890) );
  NAND3_X1 U12173 ( .A1(n15749), .A2(n15750), .A3(n15751), .ZN(n3888) );
  NAND3_X1 U12174 ( .A1(n15754), .A2(n15755), .A3(n15756), .ZN(n3886) );
  NAND3_X1 U12175 ( .A1(n15759), .A2(n15760), .A3(n15761), .ZN(n3884) );
  NAND3_X1 U12176 ( .A1(n15764), .A2(n15765), .A3(n15766), .ZN(n3882) );
  NAND3_X1 U12177 ( .A1(n15769), .A2(n15770), .A3(n15771), .ZN(n3880) );
  NAND3_X1 U12178 ( .A1(n15774), .A2(n15775), .A3(n15776), .ZN(n3878) );
  NAND3_X1 U12179 ( .A1(n15779), .A2(n15780), .A3(n15781), .ZN(n3876) );
  NAND3_X1 U12180 ( .A1(n15784), .A2(n15785), .A3(n15786), .ZN(n3874) );
  NAND3_X1 U12181 ( .A1(n15789), .A2(n15790), .A3(n15791), .ZN(n3872) );
  NAND3_X1 U12182 ( .A1(n15794), .A2(n15795), .A3(n15796), .ZN(n3870) );
  NAND3_X1 U12183 ( .A1(n15799), .A2(n15800), .A3(n15801), .ZN(n3868) );
  NAND3_X1 U12184 ( .A1(n15804), .A2(n15805), .A3(n15806), .ZN(n3866) );
  NAND3_X1 U12185 ( .A1(n15809), .A2(n15810), .A3(n15811), .ZN(n3864) );
  NAND3_X1 U12186 ( .A1(n15814), .A2(n15815), .A3(n15816), .ZN(n3862) );
  NAND3_X1 U12187 ( .A1(n15819), .A2(n15820), .A3(n15821), .ZN(n3860) );
  NAND3_X1 U12188 ( .A1(n15824), .A2(n15825), .A3(n15826), .ZN(n3858) );
  NAND3_X1 U12189 ( .A1(n15839), .A2(n14125), .A3(n15646), .ZN(n15841) );
  NAND3_X1 U12190 ( .A1(n14049), .A2(n17382), .A3(n17313), .ZN(n14186) );
  NAND3_X1 U12191 ( .A1(n15844), .A2(n15845), .A3(n15830), .ZN(n15843) );
  OAI33_X1 U12192 ( .A1(n15887), .A2(n15827), .A3(n15888), .B1(n15889), .B2(
        n15890), .B3(n15891), .ZN(n15886) );
  NAND3_X1 U12193 ( .A1(n15932), .A2(n15933), .A3(n15934), .ZN(n15892) );
  NAND3_X1 U12194 ( .A1(n15958), .A2(n15959), .A3(n15960), .ZN(n15942) );
  NAND3_X1 U12195 ( .A1(n15977), .A2(n15978), .A3(n15979), .ZN(n15961) );
  NAND3_X1 U12196 ( .A1(n15996), .A2(n15997), .A3(n15998), .ZN(n15980) );
  NAND3_X1 U12197 ( .A1(n16021), .A2(n16022), .A3(n16023), .ZN(n16005) );
  NAND3_X1 U12198 ( .A1(n16040), .A2(n16041), .A3(n16042), .ZN(n16024) );
  NAND3_X1 U12199 ( .A1(n16059), .A2(n16060), .A3(n16061), .ZN(n16043) );
  NAND3_X1 U12200 ( .A1(n16078), .A2(n16079), .A3(n16080), .ZN(n16062) );
  NAND3_X1 U12201 ( .A1(n16097), .A2(n16098), .A3(n16099), .ZN(n16081) );
  NAND3_X1 U12202 ( .A1(n16116), .A2(n16117), .A3(n16118), .ZN(n16100) );
  NAND3_X1 U12203 ( .A1(n16135), .A2(n16136), .A3(n16137), .ZN(n16119) );
  NAND3_X1 U12204 ( .A1(n16154), .A2(n16155), .A3(n16156), .ZN(n16138) );
  NAND3_X1 U12205 ( .A1(n16173), .A2(n16174), .A3(n16175), .ZN(n16157) );
  NAND3_X1 U12206 ( .A1(n16192), .A2(n16193), .A3(n16194), .ZN(n16176) );
  NAND3_X1 U12207 ( .A1(n16211), .A2(n16212), .A3(n16213), .ZN(n16195) );
  NAND3_X1 U12208 ( .A1(n16230), .A2(n16231), .A3(n16232), .ZN(n16214) );
  NAND3_X1 U12209 ( .A1(n16249), .A2(n16250), .A3(n16251), .ZN(n16233) );
  NAND3_X1 U12210 ( .A1(n16268), .A2(n16269), .A3(n16270), .ZN(n16252) );
  NAND3_X1 U12211 ( .A1(n16287), .A2(n16288), .A3(n16289), .ZN(n16271) );
  NAND3_X1 U12212 ( .A1(n16306), .A2(n16307), .A3(n16308), .ZN(n16290) );
  NAND3_X1 U12213 ( .A1(n16326), .A2(n16327), .A3(n16328), .ZN(n16310) );
  NAND3_X1 U12214 ( .A1(n16345), .A2(n16346), .A3(n16347), .ZN(n16329) );
  NAND3_X1 U12215 ( .A1(n16364), .A2(n16365), .A3(n16366), .ZN(n16348) );
  NAND3_X1 U12216 ( .A1(n16383), .A2(n16384), .A3(n16385), .ZN(n16367) );
  NAND3_X1 U12217 ( .A1(n16398), .A2(n16399), .A3(n16400), .ZN(n16387) );
  NAND3_X1 U12218 ( .A1(n16417), .A2(n16418), .A3(n16419), .ZN(n16406) );
  NAND3_X1 U12219 ( .A1(n16440), .A2(n16441), .A3(n16442), .ZN(n16424) );
  NAND3_X1 U12220 ( .A1(n16459), .A2(n16460), .A3(n16461), .ZN(n16443) );
  NAND3_X1 U12221 ( .A1(n16478), .A2(n16479), .A3(n16480), .ZN(n16462) );
  NAND3_X1 U12222 ( .A1(n16497), .A2(n16498), .A3(n16499), .ZN(n16481) );
  NAND3_X1 U12223 ( .A1(n16516), .A2(n16517), .A3(n16518), .ZN(n16500) );
  NAND3_X1 U12224 ( .A1(\pipeline/stageD/offset_jump_sign_ext [21]), .A2(
        n17384), .A3(n17328), .ZN(n16528) );
  NAND3_X1 U12225 ( .A1(n17384), .A2(n17328), .A3(n17315), .ZN(n16531) );
  NAND3_X1 U12226 ( .A1(\pipeline/stageD/offset_jump_sign_ext [24]), .A2(
        \pipeline/stageD/offset_jump_sign_ext [21]), .A3(n17328), .ZN(n16534)
         );
  NAND3_X1 U12227 ( .A1(\pipeline/stageD/offset_jump_sign_ext [31]), .A2(
        n17384), .A3(n17315), .ZN(n16539) );
  NAND3_X1 U12228 ( .A1(\pipeline/stageD/offset_jump_sign_ext [31]), .A2(
        \pipeline/stageD/offset_jump_sign_ext [21]), .A3(n17384), .ZN(n16540)
         );
  NAND3_X1 U12229 ( .A1(n16547), .A2(n16548), .A3(n16549), .ZN(n16519) );
  NAND3_X1 U12230 ( .A1(\pipeline/stageD/offset_jump_sign_ext [24]), .A2(
        n17328), .A3(n17315), .ZN(n16533) );
  NAND3_X1 U12231 ( .A1(\pipeline/stageD/offset_jump_sign_ext [31]), .A2(
        \pipeline/stageD/offset_jump_sign_ext [24]), .A3(n17315), .ZN(n16545)
         );
  NAND3_X1 U12232 ( .A1(\pipeline/stageD/offset_jump_sign_ext [24]), .A2(
        \pipeline/stageD/offset_jump_sign_ext [31]), .A3(
        \pipeline/stageD/offset_jump_sign_ext [21]), .ZN(n16546) );
  NAND3_X1 U12235 ( .A1(\pipeline/RegDst_to_WB[0] ), .A2(n17326), .A3(n17304), 
        .ZN(n16576) );
  NAND3_X1 U12236 ( .A1(\pipeline/RegDst_to_WB[1] ), .A2(n17314), .A3(n17326), 
        .ZN(n16578) );
  NAND3_X1 U12237 ( .A1(\pipeline/RegDst_to_WB[0] ), .A2(
        \pipeline/RegDst_to_WB[1] ), .A3(n17326), .ZN(n16579) );
  NAND3_X1 U12238 ( .A1(\pipeline/RegDst_to_WB[2] ), .A2(n17314), .A3(n17304), 
        .ZN(n16580) );
  NAND3_X1 U12239 ( .A1(\pipeline/RegDst_to_WB[2] ), .A2(
        \pipeline/RegDst_to_WB[0] ), .A3(n17304), .ZN(n16581) );
  NAND3_X1 U12240 ( .A1(\pipeline/RegDst_to_WB[2] ), .A2(
        \pipeline/RegDst_to_WB[1] ), .A3(n17314), .ZN(n16582) );
  NAND3_X1 U12242 ( .A1(\pipeline/RegDst_to_WB[0] ), .A2(
        \pipeline/RegDst_to_WB[2] ), .A3(\pipeline/RegDst_to_WB[1] ), .ZN(
        n16583) );
  NAND3_X1 U12244 ( .A1(n16657), .A2(n15432), .A3(n15430), .ZN(n16652) );
  XOR2_X1 U12245 ( .A(n17381), .B(n15553), .Z(n16677) );
  XOR2_X1 U12246 ( .A(n17381), .B(n15512), .Z(n15521) );
  XOR2_X1 U12247 ( .A(n17381), .B(n15474), .Z(n16666) );
  XOR2_X1 U12248 ( .A(n17381), .B(n15449), .Z(n15459) );
  XOR2_X1 U12249 ( .A(n17381), .B(n15346), .Z(n15348) );
  XOR2_X1 U12250 ( .A(n17381), .B(n15312), .Z(n16629) );
  XOR2_X1 U12251 ( .A(n17381), .B(n15285), .Z(n16626) );
  XOR2_X1 U12252 ( .A(n17381), .B(n15261), .Z(n15263) );
  XOR2_X1 U12253 ( .A(n17381), .B(n15224), .Z(n15234) );
  XOR2_X1 U12254 ( .A(n17381), .B(n15216), .Z(n16612) );
  XOR2_X1 U12255 ( .A(n17381), .B(n15202), .Z(n15204) );
  XOR2_X1 U12256 ( .A(n17381), .B(n15182), .Z(n16611) );
  NAND3_X1 U12257 ( .A1(n16789), .A2(n16790), .A3(n16791), .ZN(n16785) );
  XOR2_X1 U12258 ( .A(n17645), .B(\pipeline/Reg2_Addr_to_exe [1]), .Z(n16791)
         );
  XOR2_X1 U12259 ( .A(n17646), .B(\pipeline/Reg2_Addr_to_exe [2]), .Z(n16790)
         );
  XOR2_X1 U12261 ( .A(\pipeline/regDst_to_mem[0] ), .B(
        \pipeline/Reg1_Addr_to_exe [0]), .Z(n16809) );
  IRAM getInstr ( .ck(Clk), .Rst(n13281), .Addr({addr_to_iram[31:2], 
        \pipeline/stageF/PC_plus4/N8 , \pipeline/stageF/PC_plus4/N7 }), .Dout(
        InstrFetched) );
  TBUF_X1 \pipeline/stageD/evaluate_jump_target/targetJump_out_adder_tri[30]  ( 
        .A(\pipeline/stageD/evaluate_jump_target/N63 ), .EN(n13281), .Z(
        \pipeline/stageD/target_Jump_temp [30]) );
  TBUF_X1 \pipeline/stageD/evaluate_jump_target/targetJump_out_adder_tri[19]  ( 
        .A(\pipeline/stageD/evaluate_jump_target/N52 ), .EN(n13281), .Z(
        \pipeline/stageD/target_Jump_temp [19]) );
  TBUF_X1 \pipeline/stageD/evaluate_jump_target/targetJump_out_adder_tri[21]  ( 
        .A(\pipeline/stageD/evaluate_jump_target/N54 ), .EN(n13281), .Z(
        \pipeline/stageD/target_Jump_temp [21]) );
  TBUF_X1 \pipeline/stageD/evaluate_jump_target/targetJump_out_adder_tri[22]  ( 
        .A(\pipeline/stageD/evaluate_jump_target/N55 ), .EN(n13281), .Z(
        \pipeline/stageD/target_Jump_temp [22]) );
  NAND3_X1 U12260 ( .A1(n17314), .A2(n17326), .A3(n17304), .ZN(n16586) );
  DFF_X1 \pipeline/IFID_stage/PC_out_IFID_reg[0]  ( .D(n3879), .CK(Clk), .Q(
        \pipeline/nextPC_IFID_DEC[0] ), .QN(n17450) );
  DFF_X1 \pipeline/IFID_stage/Instr_out_IFID_reg[24]  ( .D(n3964), .CK(Clk), 
        .Q(\pipeline/stageD/offset_jump_sign_ext [24]), .QN(n17384) );
  DFF_X1 \pipeline/IFID_stage/Instr_out_IFID_reg[29]  ( .D(n3959), .CK(Clk), 
        .Q(\pipeline/inst_IFID_DEC[29] ), .QN(n17382) );
  DFF_X1 \pipeline/IFID_stage/Instr_out_IFID_reg[5]  ( .D(n3982), .CK(Clk), 
        .Q(\pipeline/stageD/offset_to_jump_temp [5]), .QN(n17350) );
  DFF_X1 \pipeline/IFID_stage/Instr_out_IFID_reg[25]  ( .D(n3963), .CK(Clk), 
        .Q(\pipeline/stageD/offset_jump_sign_ext [31]), .QN(n17328) );
  DFF_X2 \pipeline/IDEX_Stage/EXE_controls_out_IDEX_reg[0]  ( .D(
        \pipeline/IDEX_Stage/N93 ), .CK(Clk), .Q(
        \pipeline/EXE_controls_in_EXEcute [0]), .QN(n17327) );
  DFF_X1 \pipeline/MEMWB_Stage/RegDst_Addr_out_MEMWB_reg[2]  ( .D(
        \pipeline/MEMWB_Stage/N45 ), .CK(Clk), .Q(\pipeline/RegDst_to_WB[2] ), 
        .QN(n17326) );
  DFF_X1 \pipeline/IFID_stage/Instr_out_IFID_reg[22]  ( .D(n3966), .CK(Clk), 
        .Q(\pipeline/stageD/offset_jump_sign_ext [22]), .QN(n17317) );
  DFF_X1 \pipeline/IFID_stage/Instr_out_IFID_reg[21]  ( .D(n3967), .CK(Clk), 
        .Q(\pipeline/stageD/offset_jump_sign_ext [21]), .QN(n17315) );
  DFF_X1 \pipeline/IFID_stage/Instr_out_IFID_reg[27]  ( .D(n3961), .CK(Clk), 
        .Q(\pipeline/inst_IFID_DEC[27] ), .QN(n17313) );
  TBUF_X1 \DataMem/Dataout_tri[31]  ( .A(\DataMem/N2256 ), .EN(\DataMem/N0 ), 
        .Z(data_from_dram[31]) );
  TBUF_X1 \DataMem/Dataout_tri[30]  ( .A(\DataMem/N2259 ), .EN(\DataMem/N1 ), 
        .Z(data_from_dram[30]) );
  TBUF_X1 \DataMem/Dataout_tri[29]  ( .A(\DataMem/N2262 ), .EN(\DataMem/N2 ), 
        .Z(data_from_dram[29]) );
  TBUF_X1 \DataMem/Dataout_tri[28]  ( .A(\DataMem/N2265 ), .EN(\DataMem/N3 ), 
        .Z(data_from_dram[28]) );
  TBUF_X1 \DataMem/Dataout_tri[27]  ( .A(\DataMem/N2268 ), .EN(\DataMem/N4 ), 
        .Z(data_from_dram[27]) );
  TBUF_X1 \DataMem/Dataout_tri[26]  ( .A(\DataMem/N2271 ), .EN(\DataMem/N5 ), 
        .Z(data_from_dram[26]) );
  TBUF_X1 \DataMem/Dataout_tri[25]  ( .A(\DataMem/N2274 ), .EN(\DataMem/N6 ), 
        .Z(data_from_dram[25]) );
  TBUF_X1 \DataMem/Dataout_tri[24]  ( .A(\DataMem/N2277 ), .EN(\DataMem/N7 ), 
        .Z(data_from_dram[24]) );
  TBUF_X1 \DataMem/Dataout_tri[23]  ( .A(\DataMem/N2280 ), .EN(\DataMem/N8 ), 
        .Z(data_from_dram[23]) );
  TBUF_X1 \DataMem/Dataout_tri[22]  ( .A(\DataMem/N2283 ), .EN(\DataMem/N9 ), 
        .Z(data_from_dram[22]) );
  TBUF_X1 \DataMem/Dataout_tri[21]  ( .A(\DataMem/N2286 ), .EN(\DataMem/N10 ), 
        .Z(data_from_dram[21]) );
  TBUF_X1 \DataMem/Dataout_tri[20]  ( .A(\DataMem/N2289 ), .EN(\DataMem/N11 ), 
        .Z(data_from_dram[20]) );
  TBUF_X1 \DataMem/Dataout_tri[19]  ( .A(\DataMem/N2292 ), .EN(\DataMem/N12 ), 
        .Z(data_from_dram[19]) );
  TBUF_X1 \DataMem/Dataout_tri[18]  ( .A(\DataMem/N2295 ), .EN(\DataMem/N13 ), 
        .Z(data_from_dram[18]) );
  TBUF_X1 \DataMem/Dataout_tri[17]  ( .A(\DataMem/N2298 ), .EN(\DataMem/N14 ), 
        .Z(data_from_dram[17]) );
  TBUF_X1 \DataMem/Dataout_tri[16]  ( .A(\DataMem/N2301 ), .EN(\DataMem/N15 ), 
        .Z(data_from_dram[16]) );
  TBUF_X1 \DataMem/Dataout_tri[15]  ( .A(\DataMem/N2304 ), .EN(\DataMem/N16 ), 
        .Z(data_from_dram[15]) );
  TBUF_X1 \DataMem/Dataout_tri[14]  ( .A(\DataMem/N2307 ), .EN(\DataMem/N17 ), 
        .Z(data_from_dram[14]) );
  TBUF_X1 \DataMem/Dataout_tri[13]  ( .A(\DataMem/N2310 ), .EN(\DataMem/N18 ), 
        .Z(data_from_dram[13]) );
  TBUF_X1 \DataMem/Dataout_tri[12]  ( .A(\DataMem/N2313 ), .EN(\DataMem/N19 ), 
        .Z(data_from_dram[12]) );
  TBUF_X1 \DataMem/Dataout_tri[11]  ( .A(\DataMem/N2316 ), .EN(\DataMem/N20 ), 
        .Z(data_from_dram[11]) );
  TBUF_X1 \DataMem/Dataout_tri[10]  ( .A(\DataMem/N2319 ), .EN(\DataMem/N21 ), 
        .Z(data_from_dram[10]) );
  TBUF_X1 \DataMem/Dataout_tri[9]  ( .A(\DataMem/N2322 ), .EN(\DataMem/N22 ), 
        .Z(data_from_dram[9]) );
  TBUF_X1 \DataMem/Dataout_tri[8]  ( .A(\DataMem/N2325 ), .EN(\DataMem/N23 ), 
        .Z(data_from_dram[8]) );
  TBUF_X1 \DataMem/Dataout_tri[7]  ( .A(\DataMem/N2328 ), .EN(\DataMem/N24 ), 
        .Z(data_from_dram[7]) );
  TBUF_X1 \DataMem/Dataout_tri[6]  ( .A(\DataMem/N2331 ), .EN(\DataMem/N25 ), 
        .Z(data_from_dram[6]) );
  TBUF_X1 \DataMem/Dataout_tri[5]  ( .A(\DataMem/N2334 ), .EN(\DataMem/N26 ), 
        .Z(data_from_dram[5]) );
  TBUF_X1 \DataMem/Dataout_tri[4]  ( .A(\DataMem/N2337 ), .EN(\DataMem/N27 ), 
        .Z(data_from_dram[4]) );
  TBUF_X1 \DataMem/Dataout_tri[3]  ( .A(\DataMem/N2340 ), .EN(\DataMem/N28 ), 
        .Z(data_from_dram[3]) );
  TBUF_X1 \DataMem/Dataout_tri[2]  ( .A(\DataMem/N2343 ), .EN(\DataMem/N29 ), 
        .Z(data_from_dram[2]) );
  TBUF_X1 \DataMem/Dataout_tri[1]  ( .A(\DataMem/N2346 ), .EN(\DataMem/N30 ), 
        .Z(data_from_dram[1]) );
  TBUF_X1 \DataMem/Dataout_tri[0]  ( .A(\DataMem/N2349 ), .EN(\DataMem/N31 ), 
        .Z(data_from_dram[0]) );
  TBUF_X1 \pipeline/stageD/evaluate_jump_target/targetJump_out_adder_tri[31]  ( 
        .A(1'b0), .EN(n13281), .Z(\pipeline/stageD/target_Jump_temp [31]) );
  TBUF_X1 \pipeline/stageD/evaluate_jump_target/targetJump_out_adder_tri[1]  ( 
        .A(\pipeline/stageD/evaluate_jump_target/N34 ), .EN(n13281), .Z(
        \pipeline/stageD/target_Jump_temp [1]) );
  TBUF_X1 \pipeline/stageD/evaluate_jump_target/targetJump_out_adder_tri[0]  ( 
        .A(\pipeline/stageD/evaluate_jump_target/N33 ), .EN(n13281), .Z(
        \pipeline/stageD/target_Jump_temp [0]) );
  TBUF_X1 \pipeline/stageD/evaluate_jump_target/targetJump_out_adder_tri[11]  ( 
        .A(\pipeline/stageD/evaluate_jump_target/N44 ), .EN(n13281), .Z(
        \pipeline/stageD/target_Jump_temp [11]) );
  TBUF_X1 \pipeline/stageD/evaluate_jump_target/targetJump_out_adder_tri[12]  ( 
        .A(\pipeline/stageD/evaluate_jump_target/N45 ), .EN(n13281), .Z(
        \pipeline/stageD/target_Jump_temp [12]) );
  TBUF_X1 \pipeline/stageD/evaluate_jump_target/targetJump_out_adder_tri[8]  ( 
        .A(\pipeline/stageD/evaluate_jump_target/N41 ), .EN(n13281), .Z(
        \pipeline/stageD/target_Jump_temp [8]) );
  TBUF_X1 \pipeline/stageD/evaluate_jump_target/targetJump_out_adder_tri[7]  ( 
        .A(\pipeline/stageD/evaluate_jump_target/N40 ), .EN(n13281), .Z(
        \pipeline/stageD/target_Jump_temp [7]) );
  TBUF_X1 \pipeline/stageD/evaluate_jump_target/targetJump_out_adder_tri[6]  ( 
        .A(\pipeline/stageD/evaluate_jump_target/N39 ), .EN(n13281), .Z(
        \pipeline/stageD/target_Jump_temp [6]) );
  TBUF_X1 \pipeline/stageD/evaluate_jump_target/targetJump_out_adder_tri[15]  ( 
        .A(\pipeline/stageD/evaluate_jump_target/N48 ), .EN(n13281), .Z(
        \pipeline/stageD/target_Jump_temp [15]) );
  TBUF_X1 \pipeline/stageD/evaluate_jump_target/targetJump_out_adder_tri[13]  ( 
        .A(\pipeline/stageD/evaluate_jump_target/N46 ), .EN(n13281), .Z(
        \pipeline/stageD/target_Jump_temp [13]) );
  TBUF_X1 \pipeline/stageD/evaluate_jump_target/targetJump_out_adder_tri[9]  ( 
        .A(\pipeline/stageD/evaluate_jump_target/N42 ), .EN(n13281), .Z(
        \pipeline/stageD/target_Jump_temp [9]) );
  TBUF_X1 \pipeline/stageD/evaluate_jump_target/targetJump_out_adder_tri[5]  ( 
        .A(\pipeline/stageD/evaluate_jump_target/N38 ), .EN(n13281), .Z(
        \pipeline/stageD/target_Jump_temp [5]) );
  TBUF_X1 \pipeline/stageD/evaluate_jump_target/targetJump_out_adder_tri[3]  ( 
        .A(\pipeline/stageD/evaluate_jump_target/N36 ), .EN(n13281), .Z(
        \pipeline/stageD/target_Jump_temp [3]) );
  TBUF_X1 \pipeline/stageD/evaluate_jump_target/targetJump_out_adder_tri[14]  ( 
        .A(\pipeline/stageD/evaluate_jump_target/N47 ), .EN(n13281), .Z(
        \pipeline/stageD/target_Jump_temp [14]) );
  TBUF_X1 \pipeline/stageD/evaluate_jump_target/targetJump_out_adder_tri[2]  ( 
        .A(\pipeline/stageD/evaluate_jump_target/N35 ), .EN(n13281), .Z(
        \pipeline/stageD/target_Jump_temp [2]) );
  TBUF_X1 \pipeline/stageD/evaluate_jump_target/targetJump_out_adder_tri[10]  ( 
        .A(\pipeline/stageD/evaluate_jump_target/N43 ), .EN(n13281), .Z(
        \pipeline/stageD/target_Jump_temp [10]) );
  TBUF_X1 \pipeline/stageD/evaluate_jump_target/targetJump_out_adder_tri[4]  ( 
        .A(\pipeline/stageD/evaluate_jump_target/N37 ), .EN(n13281), .Z(
        \pipeline/stageD/target_Jump_temp [4]) );
  TBUF_X1 \pipeline/stageD/evaluate_jump_target/targetJump_out_adder_tri[29]  ( 
        .A(\pipeline/stageD/evaluate_jump_target/N62 ), .EN(n13281), .Z(
        \pipeline/stageD/target_Jump_temp [29]) );
  TBUF_X1 \pipeline/stageD/evaluate_jump_target/targetJump_out_adder_tri[17]  ( 
        .A(\pipeline/stageD/evaluate_jump_target/N50 ), .EN(n13281), .Z(
        \pipeline/stageD/target_Jump_temp [17]) );
  TBUF_X1 \pipeline/stageD/evaluate_jump_target/targetJump_out_adder_tri[16]  ( 
        .A(\pipeline/stageD/evaluate_jump_target/N49 ), .EN(n13281), .Z(
        \pipeline/stageD/target_Jump_temp [16]) );
  TBUF_X1 \pipeline/stageD/evaluate_jump_target/targetJump_out_adder_tri[23]  ( 
        .A(\pipeline/stageD/evaluate_jump_target/N56 ), .EN(n13281), .Z(
        \pipeline/stageD/target_Jump_temp [23]) );
  TBUF_X1 \pipeline/stageD/evaluate_jump_target/targetJump_out_adder_tri[26]  ( 
        .A(\pipeline/stageD/evaluate_jump_target/N59 ), .EN(n13281), .Z(
        \pipeline/stageD/target_Jump_temp [26]) );
  TBUF_X1 \pipeline/stageD/evaluate_jump_target/targetJump_out_adder_tri[28]  ( 
        .A(\pipeline/stageD/evaluate_jump_target/N61 ), .EN(n13281), .Z(
        \pipeline/stageD/target_Jump_temp [28]) );
  TBUF_X1 \pipeline/stageD/evaluate_jump_target/targetJump_out_adder_tri[27]  ( 
        .A(\pipeline/stageD/evaluate_jump_target/N60 ), .EN(n13281), .Z(
        \pipeline/stageD/target_Jump_temp [27]) );
  TBUF_X1 \pipeline/stageD/evaluate_jump_target/targetJump_out_adder_tri[25]  ( 
        .A(\pipeline/stageD/evaluate_jump_target/N58 ), .EN(n13281), .Z(
        \pipeline/stageD/target_Jump_temp [25]) );
  TBUF_X1 \pipeline/stageD/evaluate_jump_target/targetJump_out_adder_tri[20]  ( 
        .A(\pipeline/stageD/evaluate_jump_target/N53 ), .EN(n13281), .Z(
        \pipeline/stageD/target_Jump_temp [20]) );
  TBUF_X1 \pipeline/stageD/evaluate_jump_target/targetJump_out_adder_tri[18]  ( 
        .A(\pipeline/stageD/evaluate_jump_target/N51 ), .EN(n13281), .Z(
        \pipeline/stageD/target_Jump_temp [18]) );
  TBUF_X1 \pipeline/stageD/evaluate_jump_target/targetJump_out_adder_tri[24]  ( 
        .A(\pipeline/stageD/evaluate_jump_target/N57 ), .EN(n13281), .Z(
        \pipeline/stageD/target_Jump_temp [24]) );
  DFF_X1 \pipeline/EXMEM_stage/RegDst_Addr_out_EXMEM_reg[1]  ( .D(
        \pipeline/EXMEM_stage/N72 ), .CK(Clk), .Q(\pipeline/regDst_to_mem[1] ), 
        .QN(n17645) );
  DFF_X1 \pipeline/EXMEM_stage/RegDst_Addr_out_EXMEM_reg[2]  ( .D(
        \pipeline/EXMEM_stage/N73 ), .CK(Clk), .QN(n17646) );
  DFF_X1 \pipeline/MEMWB_Stage/RegDst_Addr_out_MEMWB_reg[0]  ( .D(
        \pipeline/MEMWB_Stage/N43 ), .CK(Clk), .Q(\pipeline/RegDst_to_WB[0] ), 
        .QN(n17314) );
  OAI21_X1 U8434 ( .B1(n13967), .B2(n17317), .A(n13969), .ZN(
        \pipeline/stageD/offset_to_jump_temp [22]) );
  OAI21_X1 U8437 ( .B1(n17349), .B2(n13967), .A(n13969), .ZN(
        \pipeline/stageD/offset_to_jump_temp [19]) );
  OAI21_X1 U8438 ( .B1(n17408), .B2(n13967), .A(n13969), .ZN(
        \pipeline/stageD/offset_to_jump_temp [18]) );
  OAI21_X1 U8439 ( .B1(n17329), .B2(n13967), .A(n13969), .ZN(
        \pipeline/stageD/offset_to_jump_temp [17]) );
  OAI21_X1 U8440 ( .B1(n17316), .B2(n13967), .A(n13969), .ZN(
        \pipeline/stageD/offset_to_jump_temp [16]) );
  OAI21_X1 U8436 ( .B1(n17407), .B2(n13967), .A(n13969), .ZN(
        \pipeline/stageD/offset_to_jump_temp [20]) );
  OAI21_X1 U8435 ( .B1(n13967), .B2(n17315), .A(n13969), .ZN(
        \pipeline/stageD/offset_to_jump_temp [21]) );
  OAI21_X1 U8433 ( .B1(n13967), .B2(n17383), .A(n13969), .ZN(
        \pipeline/stageD/offset_to_jump_temp [23]) );
  OAI21_X1 U8432 ( .B1(n13967), .B2(n17384), .A(n13969), .ZN(
        \pipeline/stageD/offset_to_jump_temp [24]) );
  OAI22_X1 U10941 ( .A1(\pipeline/regDst_to_mem[0] ), .A2(n17315), .B1(n17646), 
        .B2(\pipeline/stageD/offset_jump_sign_ext [23]), .ZN(n16575) );
  AOI221_X1 U10940 ( .B1(n17315), .B2(\pipeline/regDst_to_mem[0] ), .C1(n17646), .C2(\pipeline/stageD/offset_jump_sign_ext [23]), .A(n16575), .ZN(n16574) );
  OAI221_X1 U10937 ( .B1(\pipeline/regDst_to_mem[1] ), .B2(n17317), .C1(n17645), .C2(\pipeline/stageD/offset_jump_sign_ext [22]), .A(n16572), .ZN(n16555) );
  AOI22_X1 U10935 ( .A1(n17385), .A2(
        \pipeline/stageD/offset_jump_sign_ext [24]), .B1(n17314), .B2(
        \pipeline/stageD/offset_jump_sign_ext [21]), .ZN(n16571) );
  OAI221_X1 U10934 ( .B1(n17385), .B2(
        \pipeline/stageD/offset_jump_sign_ext [24]), .C1(n17314), .C2(
        \pipeline/stageD/offset_jump_sign_ext [21]), .A(n16571), .ZN(n16562)
         );
  NOR4_X1 U10928 ( .A1(\pipeline/Alu_Out_Addr_to_mem[19] ), .A2(
        \pipeline/Alu_Out_Addr_to_mem[18] ), .A3(
        \pipeline/Alu_Out_Addr_to_mem[20] ), .A4(
        \pipeline/Alu_Out_Addr_to_mem[21] ), .ZN(n16556) );
  NOR4_X1 U10927 ( .A1(\pipeline/Alu_Out_Addr_to_mem[25] ), .A2(
        \pipeline/Alu_Out_Addr_to_mem[24] ), .A3(
        \pipeline/Alu_Out_Addr_to_mem[23] ), .A4(
        \pipeline/Alu_Out_Addr_to_mem[22] ), .ZN(n16557) );
  NOR4_X1 U10926 ( .A1(\pipeline/Alu_Out_Addr_to_mem[13] ), .A2(
        \pipeline/Alu_Out_Addr_to_mem[11] ), .A3(
        \pipeline/Alu_Out_Addr_to_mem[10] ), .A4(
        \pipeline/Alu_Out_Addr_to_mem[12] ), .ZN(n16558) );
  NOR4_X1 U10925 ( .A1(\pipeline/Alu_Out_Addr_to_mem[14] ), .A2(
        \pipeline/Alu_Out_Addr_to_mem[15] ), .A3(
        \pipeline/Alu_Out_Addr_to_mem[17] ), .A4(
        \pipeline/Alu_Out_Addr_to_mem[16] ), .ZN(n16559) );
  NAND4_X1 U10924 ( .A1(n16556), .A2(n16557), .A3(n16558), .A4(n16559), .ZN(
        n15887) );
  NOR4_X1 U10921 ( .A1(\pipeline/Alu_Out_Addr_to_mem[0] ), .A2(
        \pipeline/Alu_Out_Addr_to_mem[2] ), .A3(
        \pipeline/Alu_Out_Addr_to_mem[1] ), .A4(
        \pipeline/Alu_Out_Addr_to_mem[3] ), .ZN(n16550) );
  NOR4_X1 U10920 ( .A1(\pipeline/Alu_Out_Addr_to_mem[8] ), .A2(
        \pipeline/Alu_Out_Addr_to_mem[7] ), .A3(
        \pipeline/Alu_Out_Addr_to_mem[6] ), .A4(
        \pipeline/Alu_Out_Addr_to_mem[9] ), .ZN(n16551) );
  NOR4_X1 U10919 ( .A1(\pipeline/Alu_Out_Addr_to_mem[31] ), .A2(
        \pipeline/Alu_Out_Addr_to_mem[4] ), .A3(
        \pipeline/Alu_Out_Addr_to_mem[5] ), .A4(
        \pipeline/Alu_Out_Addr_to_mem[30] ), .ZN(n16552) );
  NOR4_X1 U10918 ( .A1(\pipeline/Alu_Out_Addr_to_mem[26] ), .A2(
        \pipeline/Alu_Out_Addr_to_mem[27] ), .A3(
        \pipeline/Alu_Out_Addr_to_mem[28] ), .A4(
        \pipeline/Alu_Out_Addr_to_mem[29] ), .ZN(n16553) );
  NAND4_X1 U10917 ( .A1(n16550), .A2(n16551), .A3(n16552), .A4(n16553), .ZN(
        n15888) );
  AOI22_X1 U10913 ( .A1(n17137), .A2(\pipeline/RegFile_DEC_WB/RegBank[31][26] ), .B1(n17138), .B2(\pipeline/RegFile_DEC_WB/RegBank[30][26] ), .ZN(n16547) );
  AOI22_X1 U10909 ( .A1(n17130), .A2(\pipeline/RegFile_DEC_WB/RegBank[29][26] ), .B1(n17129), .B2(\pipeline/RegFile_DEC_WB/RegBank[28][26] ), .ZN(n16548) );
  AOI222_X1 U10904 ( .A1(n17135), .A2(\pipeline/RegFile_DEC_WB/RegBank[8][26] ), .B1(n17132), .B2(\pipeline/RegFile_DEC_WB/RegBank[25][26] ), .C1(n17127), 
        .C2(\pipeline/RegFile_DEC_WB/RegBank[24][26] ), .ZN(n16549) );
  AOI22_X1 U10900 ( .A1(n17143), .A2(\pipeline/RegFile_DEC_WB/RegBank[27][26] ), .B1(n17145), .B2(\pipeline/RegFile_DEC_WB/RegBank[26][26] ), .ZN(n16541) );
  AOI22_X1 U10897 ( .A1(n17146), .A2(\pipeline/RegFile_DEC_WB/RegBank[23][26] ), .B1(n17147), .B2(\pipeline/RegFile_DEC_WB/RegBank[22][26] ), .ZN(n16542) );
  AOI22_X1 U10894 ( .A1(n17148), .A2(\pipeline/RegFile_DEC_WB/RegBank[21][26] ), .B1(n17131), .B2(\pipeline/RegFile_DEC_WB/RegBank[20][26] ), .ZN(n16543) );
  AOI22_X1 U10891 ( .A1(n17128), .A2(\pipeline/RegFile_DEC_WB/RegBank[19][26] ), .B1(n17134), .B2(\pipeline/RegFile_DEC_WB/RegBank[18][26] ), .ZN(n16544) );
  NAND4_X1 U10890 ( .A1(n16541), .A2(n16542), .A3(n16543), .A4(n16544), .ZN(
        n16520) );
  AOI22_X1 U10887 ( .A1(n17141), .A2(\pipeline/RegFile_DEC_WB/RegBank[17][26] ), .B1(n17341), .B2(\pipeline/RegFile_DEC_WB/RegBank[16][26] ), .ZN(n16535) );
  AOI22_X1 U10884 ( .A1(n17388), .A2(\pipeline/RegFile_DEC_WB/RegBank[9][26] ), 
        .B1(n17139), .B2(\pipeline/RegFile_DEC_WB/RegBank[2][26] ), .ZN(n16536) );
  AOI22_X1 U10881 ( .A1(n17136), .A2(\pipeline/RegFile_DEC_WB/RegBank[12][26] ), .B1(n17389), .B2(\pipeline/RegFile_DEC_WB/RegBank[11][26] ), .ZN(n16537) );
  AOI22_X1 U10878 ( .A1(n17140), .A2(\pipeline/RegFile_DEC_WB/RegBank[14][26] ), .B1(n17390), .B2(\pipeline/RegFile_DEC_WB/RegBank[15][26] ), .ZN(n16538) );
  NAND4_X1 U10877 ( .A1(n16535), .A2(n16536), .A3(n16537), .A4(n16538), .ZN(
        n16521) );
  AOI22_X1 U10874 ( .A1(n17133), .A2(\pipeline/RegFile_DEC_WB/RegBank[13][26] ), .B1(n17392), .B2(\pipeline/RegFile_DEC_WB/RegBank[4][26] ), .ZN(n16523) );
  AOI22_X1 U10871 ( .A1(n17334), .A2(\pipeline/RegFile_DEC_WB/RegBank[10][26] ), .B1(n17144), .B2(\pipeline/RegFile_DEC_WB/RegBank[3][26] ), .ZN(n16524) );
  AOI22_X1 U10868 ( .A1(n17338), .A2(\pipeline/RegFile_DEC_WB/RegBank[6][26] ), 
        .B1(n17142), .B2(\pipeline/RegFile_DEC_WB/RegBank[7][26] ), .ZN(n16525) );
  AOI22_X1 U10865 ( .A1(n17336), .A2(\pipeline/RegFile_DEC_WB/RegBank[5][26] ), 
        .B1(n17391), .B2(\pipeline/RegFile_DEC_WB/RegBank[1][26] ), .ZN(n16526) );
  NAND4_X1 U10864 ( .A1(n16523), .A2(n16524), .A3(n16525), .A4(n16526), .ZN(
        n16522) );
  NOR4_X1 U10863 ( .A1(n16519), .A2(n16520), .A3(n16521), .A4(n16522), .ZN(
        n14893) );
  AOI22_X1 U10862 ( .A1(n15940), .A2(\pipeline/RegFile_DEC_WB/RegBank[31][25] ), .B1(n15941), .B2(\pipeline/RegFile_DEC_WB/RegBank[30][25] ), .ZN(n16516) );
  AOI22_X1 U10861 ( .A1(n15938), .A2(\pipeline/RegFile_DEC_WB/RegBank[29][25] ), .B1(n15939), .B2(\pipeline/RegFile_DEC_WB/RegBank[28][25] ), .ZN(n16517) );
  AOI222_X1 U10860 ( .A1(n15935), .A2(\pipeline/RegFile_DEC_WB/RegBank[8][25] ), .B1(n15936), .B2(\pipeline/RegFile_DEC_WB/RegBank[25][25] ), .C1(n15937), 
        .C2(\pipeline/RegFile_DEC_WB/RegBank[24][25] ), .ZN(n16518) );
  AOI22_X1 U10859 ( .A1(n15930), .A2(\pipeline/RegFile_DEC_WB/RegBank[27][25] ), .B1(n15931), .B2(\pipeline/RegFile_DEC_WB/RegBank[26][25] ), .ZN(n16512) );
  AOI22_X1 U10858 ( .A1(n15928), .A2(\pipeline/RegFile_DEC_WB/RegBank[23][25] ), .B1(n15929), .B2(\pipeline/RegFile_DEC_WB/RegBank[22][25] ), .ZN(n16513) );
  AOI22_X1 U10857 ( .A1(n15926), .A2(\pipeline/RegFile_DEC_WB/RegBank[21][25] ), .B1(n15927), .B2(\pipeline/RegFile_DEC_WB/RegBank[20][25] ), .ZN(n16514) );
  AOI22_X1 U10856 ( .A1(n15924), .A2(\pipeline/RegFile_DEC_WB/RegBank[19][25] ), .B1(n15925), .B2(\pipeline/RegFile_DEC_WB/RegBank[18][25] ), .ZN(n16515) );
  NAND4_X1 U10855 ( .A1(n16512), .A2(n16513), .A3(n16514), .A4(n16515), .ZN(
        n16501) );
  AOI22_X1 U10854 ( .A1(n15918), .A2(\pipeline/RegFile_DEC_WB/RegBank[17][25] ), .B1(n17341), .B2(\pipeline/RegFile_DEC_WB/RegBank[16][25] ), .ZN(n16508) );
  AOI22_X1 U10853 ( .A1(n17388), .A2(\pipeline/RegFile_DEC_WB/RegBank[9][25] ), 
        .B1(n15917), .B2(\pipeline/RegFile_DEC_WB/RegBank[2][25] ), .ZN(n16509) );
  AOI22_X1 U10852 ( .A1(n15914), .A2(\pipeline/RegFile_DEC_WB/RegBank[12][25] ), .B1(n17389), .B2(\pipeline/RegFile_DEC_WB/RegBank[11][25] ), .ZN(n16510) );
  AOI22_X1 U10851 ( .A1(n15912), .A2(\pipeline/RegFile_DEC_WB/RegBank[14][25] ), .B1(n17390), .B2(\pipeline/RegFile_DEC_WB/RegBank[15][25] ), .ZN(n16511) );
  NAND4_X1 U10850 ( .A1(n16508), .A2(n16509), .A3(n16510), .A4(n16511), .ZN(
        n16502) );
  AOI22_X1 U10849 ( .A1(n15906), .A2(\pipeline/RegFile_DEC_WB/RegBank[13][25] ), .B1(n17392), .B2(\pipeline/RegFile_DEC_WB/RegBank[4][25] ), .ZN(n16504) );
  AOI22_X1 U10848 ( .A1(n17334), .A2(\pipeline/RegFile_DEC_WB/RegBank[10][25] ), .B1(n15905), .B2(\pipeline/RegFile_DEC_WB/RegBank[3][25] ), .ZN(n16505) );
  AOI22_X1 U10847 ( .A1(n17338), .A2(\pipeline/RegFile_DEC_WB/RegBank[6][25] ), 
        .B1(n15903), .B2(\pipeline/RegFile_DEC_WB/RegBank[7][25] ), .ZN(n16506) );
  AOI22_X1 U10846 ( .A1(n17336), .A2(\pipeline/RegFile_DEC_WB/RegBank[5][25] ), 
        .B1(n17391), .B2(\pipeline/RegFile_DEC_WB/RegBank[1][25] ), .ZN(n16507) );
  NAND4_X1 U10845 ( .A1(n16504), .A2(n16505), .A3(n16506), .A4(n16507), .ZN(
        n16503) );
  NOR4_X1 U10844 ( .A1(n16500), .A2(n16501), .A3(n16502), .A4(n16503), .ZN(
        n14895) );
  AOI22_X1 U10843 ( .A1(n17137), .A2(\pipeline/RegFile_DEC_WB/RegBank[31][24] ), .B1(n17138), .B2(\pipeline/RegFile_DEC_WB/RegBank[30][24] ), .ZN(n16497) );
  AOI22_X1 U10842 ( .A1(n17130), .A2(\pipeline/RegFile_DEC_WB/RegBank[29][24] ), .B1(n17129), .B2(\pipeline/RegFile_DEC_WB/RegBank[28][24] ), .ZN(n16498) );
  AOI222_X1 U10841 ( .A1(n17135), .A2(\pipeline/RegFile_DEC_WB/RegBank[8][24] ), .B1(n17132), .B2(\pipeline/RegFile_DEC_WB/RegBank[25][24] ), .C1(n17127), 
        .C2(\pipeline/RegFile_DEC_WB/RegBank[24][24] ), .ZN(n16499) );
  AOI22_X1 U10840 ( .A1(n17143), .A2(\pipeline/RegFile_DEC_WB/RegBank[27][24] ), .B1(n17145), .B2(\pipeline/RegFile_DEC_WB/RegBank[26][24] ), .ZN(n16493) );
  AOI22_X1 U10839 ( .A1(n17146), .A2(\pipeline/RegFile_DEC_WB/RegBank[23][24] ), .B1(n17147), .B2(\pipeline/RegFile_DEC_WB/RegBank[22][24] ), .ZN(n16494) );
  AOI22_X1 U10838 ( .A1(n17148), .A2(\pipeline/RegFile_DEC_WB/RegBank[21][24] ), .B1(n17131), .B2(\pipeline/RegFile_DEC_WB/RegBank[20][24] ), .ZN(n16495) );
  AOI22_X1 U10837 ( .A1(n17128), .A2(\pipeline/RegFile_DEC_WB/RegBank[19][24] ), .B1(n17134), .B2(\pipeline/RegFile_DEC_WB/RegBank[18][24] ), .ZN(n16496) );
  NAND4_X1 U10836 ( .A1(n16493), .A2(n16494), .A3(n16495), .A4(n16496), .ZN(
        n16482) );
  AOI22_X1 U10835 ( .A1(n17141), .A2(\pipeline/RegFile_DEC_WB/RegBank[17][24] ), .B1(n17341), .B2(\pipeline/RegFile_DEC_WB/RegBank[16][24] ), .ZN(n16489) );
  AOI22_X1 U10834 ( .A1(n17388), .A2(\pipeline/RegFile_DEC_WB/RegBank[9][24] ), 
        .B1(n17139), .B2(\pipeline/RegFile_DEC_WB/RegBank[2][24] ), .ZN(n16490) );
  AOI22_X1 U10833 ( .A1(n17136), .A2(\pipeline/RegFile_DEC_WB/RegBank[12][24] ), .B1(n17389), .B2(\pipeline/RegFile_DEC_WB/RegBank[11][24] ), .ZN(n16491) );
  AOI22_X1 U10832 ( .A1(n17140), .A2(\pipeline/RegFile_DEC_WB/RegBank[14][24] ), .B1(n17390), .B2(\pipeline/RegFile_DEC_WB/RegBank[15][24] ), .ZN(n16492) );
  NAND4_X1 U10831 ( .A1(n16489), .A2(n16490), .A3(n16491), .A4(n16492), .ZN(
        n16483) );
  AOI22_X1 U10830 ( .A1(n17133), .A2(\pipeline/RegFile_DEC_WB/RegBank[13][24] ), .B1(n17392), .B2(\pipeline/RegFile_DEC_WB/RegBank[4][24] ), .ZN(n16485) );
  AOI22_X1 U10829 ( .A1(n17334), .A2(\pipeline/RegFile_DEC_WB/RegBank[10][24] ), .B1(n17144), .B2(\pipeline/RegFile_DEC_WB/RegBank[3][24] ), .ZN(n16486) );
  AOI22_X1 U10828 ( .A1(n17338), .A2(\pipeline/RegFile_DEC_WB/RegBank[6][24] ), 
        .B1(n17142), .B2(\pipeline/RegFile_DEC_WB/RegBank[7][24] ), .ZN(n16487) );
  AOI22_X1 U10827 ( .A1(n17336), .A2(\pipeline/RegFile_DEC_WB/RegBank[5][24] ), 
        .B1(n17391), .B2(\pipeline/RegFile_DEC_WB/RegBank[1][24] ), .ZN(n16488) );
  NAND4_X1 U10826 ( .A1(n16485), .A2(n16486), .A3(n16487), .A4(n16488), .ZN(
        n16484) );
  NOR4_X1 U10825 ( .A1(n16481), .A2(n16482), .A3(n16483), .A4(n16484), .ZN(
        n14897) );
  AOI22_X1 U10824 ( .A1(n17137), .A2(\pipeline/RegFile_DEC_WB/RegBank[31][23] ), .B1(n17138), .B2(\pipeline/RegFile_DEC_WB/RegBank[30][23] ), .ZN(n16478) );
  AOI22_X1 U10823 ( .A1(n17130), .A2(\pipeline/RegFile_DEC_WB/RegBank[29][23] ), .B1(n17129), .B2(\pipeline/RegFile_DEC_WB/RegBank[28][23] ), .ZN(n16479) );
  AOI222_X1 U10822 ( .A1(n17135), .A2(\pipeline/RegFile_DEC_WB/RegBank[8][23] ), .B1(n17132), .B2(\pipeline/RegFile_DEC_WB/RegBank[25][23] ), .C1(n17127), 
        .C2(\pipeline/RegFile_DEC_WB/RegBank[24][23] ), .ZN(n16480) );
  AOI22_X1 U10821 ( .A1(n17143), .A2(\pipeline/RegFile_DEC_WB/RegBank[27][23] ), .B1(n17145), .B2(\pipeline/RegFile_DEC_WB/RegBank[26][23] ), .ZN(n16474) );
  AOI22_X1 U10820 ( .A1(n17146), .A2(\pipeline/RegFile_DEC_WB/RegBank[23][23] ), .B1(n17147), .B2(\pipeline/RegFile_DEC_WB/RegBank[22][23] ), .ZN(n16475) );
  AOI22_X1 U10819 ( .A1(n17148), .A2(\pipeline/RegFile_DEC_WB/RegBank[21][23] ), .B1(n17131), .B2(\pipeline/RegFile_DEC_WB/RegBank[20][23] ), .ZN(n16476) );
  AOI22_X1 U10818 ( .A1(n17128), .A2(\pipeline/RegFile_DEC_WB/RegBank[19][23] ), .B1(n17134), .B2(\pipeline/RegFile_DEC_WB/RegBank[18][23] ), .ZN(n16477) );
  NAND4_X1 U10817 ( .A1(n16474), .A2(n16475), .A3(n16476), .A4(n16477), .ZN(
        n16463) );
  AOI22_X1 U10816 ( .A1(n17141), .A2(\pipeline/RegFile_DEC_WB/RegBank[17][23] ), .B1(n17341), .B2(\pipeline/RegFile_DEC_WB/RegBank[16][23] ), .ZN(n16470) );
  AOI22_X1 U10815 ( .A1(n17388), .A2(\pipeline/RegFile_DEC_WB/RegBank[9][23] ), 
        .B1(n17139), .B2(\pipeline/RegFile_DEC_WB/RegBank[2][23] ), .ZN(n16471) );
  AOI22_X1 U10814 ( .A1(n17136), .A2(\pipeline/RegFile_DEC_WB/RegBank[12][23] ), .B1(n17389), .B2(\pipeline/RegFile_DEC_WB/RegBank[11][23] ), .ZN(n16472) );
  AOI22_X1 U10813 ( .A1(n17140), .A2(\pipeline/RegFile_DEC_WB/RegBank[14][23] ), .B1(n17390), .B2(\pipeline/RegFile_DEC_WB/RegBank[15][23] ), .ZN(n16473) );
  NAND4_X1 U10812 ( .A1(n16470), .A2(n16471), .A3(n16472), .A4(n16473), .ZN(
        n16464) );
  AOI22_X1 U10811 ( .A1(n17133), .A2(\pipeline/RegFile_DEC_WB/RegBank[13][23] ), .B1(n17392), .B2(\pipeline/RegFile_DEC_WB/RegBank[4][23] ), .ZN(n16466) );
  AOI22_X1 U10810 ( .A1(n17334), .A2(\pipeline/RegFile_DEC_WB/RegBank[10][23] ), .B1(n17144), .B2(\pipeline/RegFile_DEC_WB/RegBank[3][23] ), .ZN(n16467) );
  AOI22_X1 U10809 ( .A1(n17338), .A2(\pipeline/RegFile_DEC_WB/RegBank[6][23] ), 
        .B1(n17142), .B2(\pipeline/RegFile_DEC_WB/RegBank[7][23] ), .ZN(n16468) );
  AOI22_X1 U10808 ( .A1(n17336), .A2(\pipeline/RegFile_DEC_WB/RegBank[5][23] ), 
        .B1(n17391), .B2(\pipeline/RegFile_DEC_WB/RegBank[1][23] ), .ZN(n16469) );
  NAND4_X1 U10807 ( .A1(n16466), .A2(n16467), .A3(n16468), .A4(n16469), .ZN(
        n16465) );
  NOR4_X1 U10806 ( .A1(n16462), .A2(n16463), .A3(n16464), .A4(n16465), .ZN(
        n14899) );
  NAND4_X1 U10805 ( .A1(n14893), .A2(n14895), .A3(n14897), .A4(n14899), .ZN(
        n15889) );
  AOI22_X1 U10804 ( .A1(n17137), .A2(\pipeline/RegFile_DEC_WB/RegBank[31][6] ), 
        .B1(n17138), .B2(\pipeline/RegFile_DEC_WB/RegBank[30][6] ), .ZN(n16459) );
  AOI22_X1 U10803 ( .A1(n17130), .A2(\pipeline/RegFile_DEC_WB/RegBank[29][6] ), 
        .B1(n17129), .B2(\pipeline/RegFile_DEC_WB/RegBank[28][6] ), .ZN(n16460) );
  AOI222_X1 U10802 ( .A1(n17135), .A2(\pipeline/RegFile_DEC_WB/RegBank[8][6] ), 
        .B1(n17132), .B2(\pipeline/RegFile_DEC_WB/RegBank[25][6] ), .C1(n17127), .C2(\pipeline/RegFile_DEC_WB/RegBank[24][6] ), .ZN(n16461) );
  AOI22_X1 U10801 ( .A1(n17143), .A2(\pipeline/RegFile_DEC_WB/RegBank[27][6] ), 
        .B1(n17145), .B2(\pipeline/RegFile_DEC_WB/RegBank[26][6] ), .ZN(n16455) );
  AOI22_X1 U10800 ( .A1(n17146), .A2(\pipeline/RegFile_DEC_WB/RegBank[23][6] ), 
        .B1(n17147), .B2(\pipeline/RegFile_DEC_WB/RegBank[22][6] ), .ZN(n16456) );
  AOI22_X1 U10799 ( .A1(n17148), .A2(\pipeline/RegFile_DEC_WB/RegBank[21][6] ), 
        .B1(n17131), .B2(\pipeline/RegFile_DEC_WB/RegBank[20][6] ), .ZN(n16457) );
  AOI22_X1 U10798 ( .A1(n17128), .A2(\pipeline/RegFile_DEC_WB/RegBank[19][6] ), 
        .B1(n17134), .B2(\pipeline/RegFile_DEC_WB/RegBank[18][6] ), .ZN(n16458) );
  NAND4_X1 U10797 ( .A1(n16455), .A2(n16456), .A3(n16457), .A4(n16458), .ZN(
        n16444) );
  AOI22_X1 U10796 ( .A1(n17141), .A2(\pipeline/RegFile_DEC_WB/RegBank[17][6] ), 
        .B1(n17342), .B2(\pipeline/RegFile_DEC_WB/RegBank[16][6] ), .ZN(n16451) );
  AOI22_X1 U10795 ( .A1(n17388), .A2(\pipeline/RegFile_DEC_WB/RegBank[9][6] ), 
        .B1(n17139), .B2(\pipeline/RegFile_DEC_WB/RegBank[2][6] ), .ZN(n16452)
         );
  AOI22_X1 U10794 ( .A1(n17136), .A2(\pipeline/RegFile_DEC_WB/RegBank[12][6] ), 
        .B1(n17389), .B2(\pipeline/RegFile_DEC_WB/RegBank[11][6] ), .ZN(n16453) );
  AOI22_X1 U10793 ( .A1(n17140), .A2(\pipeline/RegFile_DEC_WB/RegBank[14][6] ), 
        .B1(n17390), .B2(\pipeline/RegFile_DEC_WB/RegBank[15][6] ), .ZN(n16454) );
  NAND4_X1 U10792 ( .A1(n16451), .A2(n16452), .A3(n16453), .A4(n16454), .ZN(
        n16445) );
  AOI22_X1 U10791 ( .A1(n17133), .A2(\pipeline/RegFile_DEC_WB/RegBank[13][6] ), 
        .B1(n17392), .B2(\pipeline/RegFile_DEC_WB/RegBank[4][6] ), .ZN(n16447)
         );
  AOI22_X1 U10790 ( .A1(n17335), .A2(\pipeline/RegFile_DEC_WB/RegBank[10][6] ), 
        .B1(n17144), .B2(\pipeline/RegFile_DEC_WB/RegBank[3][6] ), .ZN(n16448)
         );
  AOI22_X1 U10789 ( .A1(n17339), .A2(\pipeline/RegFile_DEC_WB/RegBank[6][6] ), 
        .B1(n17142), .B2(\pipeline/RegFile_DEC_WB/RegBank[7][6] ), .ZN(n16449)
         );
  AOI22_X1 U10788 ( .A1(n17337), .A2(\pipeline/RegFile_DEC_WB/RegBank[5][6] ), 
        .B1(n17391), .B2(\pipeline/RegFile_DEC_WB/RegBank[1][6] ), .ZN(n16450)
         );
  NAND4_X1 U10787 ( .A1(n16447), .A2(n16448), .A3(n16449), .A4(n16450), .ZN(
        n16446) );
  NOR4_X1 U10786 ( .A1(n16443), .A2(n16444), .A3(n16445), .A4(n16446), .ZN(
        n14933) );
  AOI22_X1 U10785 ( .A1(n15940), .A2(\pipeline/RegFile_DEC_WB/RegBank[31][5] ), 
        .B1(n15941), .B2(\pipeline/RegFile_DEC_WB/RegBank[30][5] ), .ZN(n16440) );
  AOI22_X1 U10784 ( .A1(n15938), .A2(\pipeline/RegFile_DEC_WB/RegBank[29][5] ), 
        .B1(n15939), .B2(\pipeline/RegFile_DEC_WB/RegBank[28][5] ), .ZN(n16441) );
  AOI222_X1 U10783 ( .A1(n15935), .A2(\pipeline/RegFile_DEC_WB/RegBank[8][5] ), 
        .B1(n15936), .B2(\pipeline/RegFile_DEC_WB/RegBank[25][5] ), .C1(n15937), .C2(\pipeline/RegFile_DEC_WB/RegBank[24][5] ), .ZN(n16442) );
  AOI22_X1 U10782 ( .A1(n15930), .A2(\pipeline/RegFile_DEC_WB/RegBank[27][5] ), 
        .B1(n15931), .B2(\pipeline/RegFile_DEC_WB/RegBank[26][5] ), .ZN(n16436) );
  AOI22_X1 U10781 ( .A1(n15928), .A2(\pipeline/RegFile_DEC_WB/RegBank[23][5] ), 
        .B1(n15929), .B2(\pipeline/RegFile_DEC_WB/RegBank[22][5] ), .ZN(n16437) );
  AOI22_X1 U10780 ( .A1(n15926), .A2(\pipeline/RegFile_DEC_WB/RegBank[21][5] ), 
        .B1(n15927), .B2(\pipeline/RegFile_DEC_WB/RegBank[20][5] ), .ZN(n16438) );
  AOI22_X1 U10779 ( .A1(n15924), .A2(\pipeline/RegFile_DEC_WB/RegBank[19][5] ), 
        .B1(n15925), .B2(\pipeline/RegFile_DEC_WB/RegBank[18][5] ), .ZN(n16439) );
  NAND4_X1 U10778 ( .A1(n16436), .A2(n16437), .A3(n16438), .A4(n16439), .ZN(
        n16425) );
  AOI22_X1 U10777 ( .A1(n15918), .A2(\pipeline/RegFile_DEC_WB/RegBank[17][5] ), 
        .B1(n17342), .B2(\pipeline/RegFile_DEC_WB/RegBank[16][5] ), .ZN(n16432) );
  AOI22_X1 U10776 ( .A1(n17388), .A2(\pipeline/RegFile_DEC_WB/RegBank[9][5] ), 
        .B1(n15917), .B2(\pipeline/RegFile_DEC_WB/RegBank[2][5] ), .ZN(n16433)
         );
  AOI22_X1 U10775 ( .A1(n15914), .A2(\pipeline/RegFile_DEC_WB/RegBank[12][5] ), 
        .B1(n17389), .B2(\pipeline/RegFile_DEC_WB/RegBank[11][5] ), .ZN(n16434) );
  AOI22_X1 U10774 ( .A1(n15912), .A2(\pipeline/RegFile_DEC_WB/RegBank[14][5] ), 
        .B1(n17390), .B2(\pipeline/RegFile_DEC_WB/RegBank[15][5] ), .ZN(n16435) );
  NAND4_X1 U10773 ( .A1(n16432), .A2(n16433), .A3(n16434), .A4(n16435), .ZN(
        n16426) );
  AOI22_X1 U10772 ( .A1(n15906), .A2(\pipeline/RegFile_DEC_WB/RegBank[13][5] ), 
        .B1(n17392), .B2(\pipeline/RegFile_DEC_WB/RegBank[4][5] ), .ZN(n16428)
         );
  AOI22_X1 U10771 ( .A1(n17335), .A2(\pipeline/RegFile_DEC_WB/RegBank[10][5] ), 
        .B1(n15905), .B2(\pipeline/RegFile_DEC_WB/RegBank[3][5] ), .ZN(n16429)
         );
  AOI22_X1 U10770 ( .A1(n17339), .A2(\pipeline/RegFile_DEC_WB/RegBank[6][5] ), 
        .B1(n15903), .B2(\pipeline/RegFile_DEC_WB/RegBank[7][5] ), .ZN(n16430)
         );
  AOI22_X1 U10769 ( .A1(n17337), .A2(\pipeline/RegFile_DEC_WB/RegBank[5][5] ), 
        .B1(n17391), .B2(\pipeline/RegFile_DEC_WB/RegBank[1][5] ), .ZN(n16431)
         );
  NAND4_X1 U10768 ( .A1(n16428), .A2(n16429), .A3(n16430), .A4(n16431), .ZN(
        n16427) );
  NOR4_X1 U10767 ( .A1(n16424), .A2(n16425), .A3(n16426), .A4(n16427), .ZN(
        n14935) );
  AOI22_X1 U10765 ( .A1(n15930), .A2(\pipeline/RegFile_DEC_WB/RegBank[27][0] ), 
        .B1(n15931), .B2(\pipeline/RegFile_DEC_WB/RegBank[26][0] ), .ZN(n16420) );
  AOI22_X1 U10764 ( .A1(n15928), .A2(\pipeline/RegFile_DEC_WB/RegBank[23][0] ), 
        .B1(n15929), .B2(\pipeline/RegFile_DEC_WB/RegBank[22][0] ), .ZN(n16421) );
  AOI22_X1 U10763 ( .A1(n15926), .A2(\pipeline/RegFile_DEC_WB/RegBank[21][0] ), 
        .B1(n15927), .B2(\pipeline/RegFile_DEC_WB/RegBank[20][0] ), .ZN(n16422) );
  AOI22_X1 U10762 ( .A1(n15924), .A2(\pipeline/RegFile_DEC_WB/RegBank[19][0] ), 
        .B1(n15925), .B2(\pipeline/RegFile_DEC_WB/RegBank[18][0] ), .ZN(n16423) );
  NAND4_X1 U10761 ( .A1(n16420), .A2(n16421), .A3(n16422), .A4(n16423), .ZN(
        n16405) );
  AOI22_X1 U10760 ( .A1(n15940), .A2(\pipeline/RegFile_DEC_WB/RegBank[31][0] ), 
        .B1(n15941), .B2(\pipeline/RegFile_DEC_WB/RegBank[30][0] ), .ZN(n16417) );
  AOI22_X1 U10759 ( .A1(n15938), .A2(\pipeline/RegFile_DEC_WB/RegBank[29][0] ), 
        .B1(n15939), .B2(\pipeline/RegFile_DEC_WB/RegBank[28][0] ), .ZN(n16418) );
  AOI222_X1 U10758 ( .A1(n15935), .A2(\pipeline/RegFile_DEC_WB/RegBank[8][0] ), 
        .B1(n15936), .B2(\pipeline/RegFile_DEC_WB/RegBank[25][0] ), .C1(n15937), .C2(\pipeline/RegFile_DEC_WB/RegBank[24][0] ), .ZN(n16419) );
  AOI22_X1 U10757 ( .A1(n15906), .A2(\pipeline/RegFile_DEC_WB/RegBank[13][0] ), 
        .B1(n17392), .B2(\pipeline/RegFile_DEC_WB/RegBank[4][0] ), .ZN(n16413)
         );
  AOI22_X1 U10756 ( .A1(n17335), .A2(\pipeline/RegFile_DEC_WB/RegBank[10][0] ), 
        .B1(n15905), .B2(\pipeline/RegFile_DEC_WB/RegBank[3][0] ), .ZN(n16414)
         );
  AOI22_X1 U10755 ( .A1(n17339), .A2(\pipeline/RegFile_DEC_WB/RegBank[6][0] ), 
        .B1(n15903), .B2(\pipeline/RegFile_DEC_WB/RegBank[7][0] ), .ZN(n16415)
         );
  AOI22_X1 U10754 ( .A1(n17337), .A2(\pipeline/RegFile_DEC_WB/RegBank[5][0] ), 
        .B1(n17391), .B2(\pipeline/RegFile_DEC_WB/RegBank[1][0] ), .ZN(n16416)
         );
  NAND4_X1 U10753 ( .A1(n16413), .A2(n16414), .A3(n16415), .A4(n16416), .ZN(
        n16407) );
  AOI22_X1 U10752 ( .A1(n15918), .A2(\pipeline/RegFile_DEC_WB/RegBank[17][0] ), 
        .B1(n17342), .B2(\pipeline/RegFile_DEC_WB/RegBank[16][0] ), .ZN(n16409) );
  AOI22_X1 U10751 ( .A1(n17388), .A2(\pipeline/RegFile_DEC_WB/RegBank[9][0] ), 
        .B1(n15917), .B2(\pipeline/RegFile_DEC_WB/RegBank[2][0] ), .ZN(n16410)
         );
  AOI22_X1 U10750 ( .A1(n15914), .A2(\pipeline/RegFile_DEC_WB/RegBank[12][0] ), 
        .B1(n17389), .B2(\pipeline/RegFile_DEC_WB/RegBank[11][0] ), .ZN(n16411) );
  AOI22_X1 U10749 ( .A1(n15912), .A2(\pipeline/RegFile_DEC_WB/RegBank[14][0] ), 
        .B1(n17390), .B2(\pipeline/RegFile_DEC_WB/RegBank[15][0] ), .ZN(n16412) );
  NAND4_X1 U10748 ( .A1(n16409), .A2(n16410), .A3(n16411), .A4(n16412), .ZN(
        n16408) );
  NOR4_X1 U10747 ( .A1(n16405), .A2(n16406), .A3(n16407), .A4(n16408), .ZN(
        n14945) );
  AOI22_X1 U10745 ( .A1(n17143), .A2(\pipeline/RegFile_DEC_WB/RegBank[27][31] ), .B1(n17145), .B2(\pipeline/RegFile_DEC_WB/RegBank[26][31] ), .ZN(n16401) );
  AOI22_X1 U10744 ( .A1(n17146), .A2(\pipeline/RegFile_DEC_WB/RegBank[23][31] ), .B1(n17147), .B2(\pipeline/RegFile_DEC_WB/RegBank[22][31] ), .ZN(n16402) );
  AOI22_X1 U10743 ( .A1(n17148), .A2(\pipeline/RegFile_DEC_WB/RegBank[21][31] ), .B1(n17131), .B2(\pipeline/RegFile_DEC_WB/RegBank[20][31] ), .ZN(n16403) );
  AOI22_X1 U10742 ( .A1(n17128), .A2(\pipeline/RegFile_DEC_WB/RegBank[19][31] ), .B1(n17134), .B2(\pipeline/RegFile_DEC_WB/RegBank[18][31] ), .ZN(n16404) );
  NAND4_X1 U10741 ( .A1(n16401), .A2(n16402), .A3(n16403), .A4(n16404), .ZN(
        n16386) );
  AOI22_X1 U10740 ( .A1(n17137), .A2(\pipeline/RegFile_DEC_WB/RegBank[31][31] ), .B1(n17138), .B2(\pipeline/RegFile_DEC_WB/RegBank[30][31] ), .ZN(n16398) );
  AOI22_X1 U10739 ( .A1(n17130), .A2(\pipeline/RegFile_DEC_WB/RegBank[29][31] ), .B1(n17129), .B2(\pipeline/RegFile_DEC_WB/RegBank[28][31] ), .ZN(n16399) );
  AOI222_X1 U10738 ( .A1(n17135), .A2(\pipeline/RegFile_DEC_WB/RegBank[8][31] ), .B1(n17132), .B2(\pipeline/RegFile_DEC_WB/RegBank[25][31] ), .C1(n17127), 
        .C2(\pipeline/RegFile_DEC_WB/RegBank[24][31] ), .ZN(n16400) );
  AOI22_X1 U10737 ( .A1(n17133), .A2(\pipeline/RegFile_DEC_WB/RegBank[13][31] ), .B1(n15907), .B2(\pipeline/RegFile_DEC_WB/RegBank[4][31] ), .ZN(n16394) );
  AOI22_X1 U10736 ( .A1(n17335), .A2(\pipeline/RegFile_DEC_WB/RegBank[10][31] ), .B1(n17144), .B2(\pipeline/RegFile_DEC_WB/RegBank[3][31] ), .ZN(n16395) );
  AOI22_X1 U10735 ( .A1(n17339), .A2(\pipeline/RegFile_DEC_WB/RegBank[6][31] ), 
        .B1(n17142), .B2(\pipeline/RegFile_DEC_WB/RegBank[7][31] ), .ZN(n16396) );
  AOI22_X1 U10734 ( .A1(n17337), .A2(\pipeline/RegFile_DEC_WB/RegBank[5][31] ), 
        .B1(n15901), .B2(\pipeline/RegFile_DEC_WB/RegBank[1][31] ), .ZN(n16397) );
  NAND4_X1 U10733 ( .A1(n16394), .A2(n16395), .A3(n16396), .A4(n16397), .ZN(
        n16388) );
  AOI22_X1 U10732 ( .A1(n17141), .A2(\pipeline/RegFile_DEC_WB/RegBank[17][31] ), .B1(n17342), .B2(\pipeline/RegFile_DEC_WB/RegBank[16][31] ), .ZN(n16390) );
  AOI22_X1 U10731 ( .A1(n15916), .A2(\pipeline/RegFile_DEC_WB/RegBank[9][31] ), 
        .B1(n17139), .B2(\pipeline/RegFile_DEC_WB/RegBank[2][31] ), .ZN(n16391) );
  AOI22_X1 U10730 ( .A1(n17136), .A2(\pipeline/RegFile_DEC_WB/RegBank[12][31] ), .B1(n15915), .B2(\pipeline/RegFile_DEC_WB/RegBank[11][31] ), .ZN(n16392) );
  AOI22_X1 U10729 ( .A1(n17140), .A2(\pipeline/RegFile_DEC_WB/RegBank[14][31] ), .B1(n15913), .B2(\pipeline/RegFile_DEC_WB/RegBank[15][31] ), .ZN(n16393) );
  NAND4_X1 U10728 ( .A1(n16390), .A2(n16391), .A3(n16392), .A4(n16393), .ZN(
        n16389) );
  NOR4_X1 U10727 ( .A1(n16386), .A2(n16387), .A3(n16388), .A4(n16389), .ZN(
        n14883) );
  AOI22_X1 U10725 ( .A1(n17137), .A2(\pipeline/RegFile_DEC_WB/RegBank[31][4] ), 
        .B1(n17138), .B2(\pipeline/RegFile_DEC_WB/RegBank[30][4] ), .ZN(n16383) );
  AOI22_X1 U10724 ( .A1(n17130), .A2(\pipeline/RegFile_DEC_WB/RegBank[29][4] ), 
        .B1(n17129), .B2(\pipeline/RegFile_DEC_WB/RegBank[28][4] ), .ZN(n16384) );
  AOI222_X1 U10723 ( .A1(n17135), .A2(\pipeline/RegFile_DEC_WB/RegBank[8][4] ), 
        .B1(n17132), .B2(\pipeline/RegFile_DEC_WB/RegBank[25][4] ), .C1(n17127), .C2(\pipeline/RegFile_DEC_WB/RegBank[24][4] ), .ZN(n16385) );
  AOI22_X1 U10722 ( .A1(n17143), .A2(\pipeline/RegFile_DEC_WB/RegBank[27][4] ), 
        .B1(n17145), .B2(\pipeline/RegFile_DEC_WB/RegBank[26][4] ), .ZN(n16379) );
  AOI22_X1 U10721 ( .A1(n17146), .A2(\pipeline/RegFile_DEC_WB/RegBank[23][4] ), 
        .B1(n17147), .B2(\pipeline/RegFile_DEC_WB/RegBank[22][4] ), .ZN(n16380) );
  AOI22_X1 U10720 ( .A1(n17148), .A2(\pipeline/RegFile_DEC_WB/RegBank[21][4] ), 
        .B1(n17131), .B2(\pipeline/RegFile_DEC_WB/RegBank[20][4] ), .ZN(n16381) );
  AOI22_X1 U10719 ( .A1(n17128), .A2(\pipeline/RegFile_DEC_WB/RegBank[19][4] ), 
        .B1(n17134), .B2(\pipeline/RegFile_DEC_WB/RegBank[18][4] ), .ZN(n16382) );
  NAND4_X1 U10718 ( .A1(n16379), .A2(n16380), .A3(n16381), .A4(n16382), .ZN(
        n16368) );
  AOI22_X1 U10717 ( .A1(n17141), .A2(\pipeline/RegFile_DEC_WB/RegBank[17][4] ), 
        .B1(n17342), .B2(\pipeline/RegFile_DEC_WB/RegBank[16][4] ), .ZN(n16375) );
  AOI22_X1 U10716 ( .A1(n15916), .A2(\pipeline/RegFile_DEC_WB/RegBank[9][4] ), 
        .B1(n17139), .B2(\pipeline/RegFile_DEC_WB/RegBank[2][4] ), .ZN(n16376)
         );
  AOI22_X1 U10715 ( .A1(n17136), .A2(\pipeline/RegFile_DEC_WB/RegBank[12][4] ), 
        .B1(n15915), .B2(\pipeline/RegFile_DEC_WB/RegBank[11][4] ), .ZN(n16377) );
  AOI22_X1 U10714 ( .A1(n17140), .A2(\pipeline/RegFile_DEC_WB/RegBank[14][4] ), 
        .B1(n15913), .B2(\pipeline/RegFile_DEC_WB/RegBank[15][4] ), .ZN(n16378) );
  NAND4_X1 U10713 ( .A1(n16375), .A2(n16376), .A3(n16377), .A4(n16378), .ZN(
        n16369) );
  AOI22_X1 U10712 ( .A1(n17133), .A2(\pipeline/RegFile_DEC_WB/RegBank[13][4] ), 
        .B1(n15907), .B2(\pipeline/RegFile_DEC_WB/RegBank[4][4] ), .ZN(n16371)
         );
  AOI22_X1 U10711 ( .A1(n17335), .A2(\pipeline/RegFile_DEC_WB/RegBank[10][4] ), 
        .B1(n17144), .B2(\pipeline/RegFile_DEC_WB/RegBank[3][4] ), .ZN(n16372)
         );
  AOI22_X1 U10710 ( .A1(n17339), .A2(\pipeline/RegFile_DEC_WB/RegBank[6][4] ), 
        .B1(n17142), .B2(\pipeline/RegFile_DEC_WB/RegBank[7][4] ), .ZN(n16373)
         );
  AOI22_X1 U10709 ( .A1(n17337), .A2(\pipeline/RegFile_DEC_WB/RegBank[5][4] ), 
        .B1(n15901), .B2(\pipeline/RegFile_DEC_WB/RegBank[1][4] ), .ZN(n16374)
         );
  NAND4_X1 U10708 ( .A1(n16371), .A2(n16372), .A3(n16373), .A4(n16374), .ZN(
        n16370) );
  NOR4_X1 U10707 ( .A1(n16367), .A2(n16368), .A3(n16369), .A4(n16370), .ZN(
        n14937) );
  AOI22_X1 U10706 ( .A1(n17137), .A2(\pipeline/RegFile_DEC_WB/RegBank[31][3] ), 
        .B1(n17138), .B2(\pipeline/RegFile_DEC_WB/RegBank[30][3] ), .ZN(n16364) );
  AOI22_X1 U10705 ( .A1(n17130), .A2(\pipeline/RegFile_DEC_WB/RegBank[29][3] ), 
        .B1(n17129), .B2(\pipeline/RegFile_DEC_WB/RegBank[28][3] ), .ZN(n16365) );
  AOI222_X1 U10704 ( .A1(n17135), .A2(\pipeline/RegFile_DEC_WB/RegBank[8][3] ), 
        .B1(n17132), .B2(\pipeline/RegFile_DEC_WB/RegBank[25][3] ), .C1(n17127), .C2(\pipeline/RegFile_DEC_WB/RegBank[24][3] ), .ZN(n16366) );
  AOI22_X1 U10703 ( .A1(n17143), .A2(\pipeline/RegFile_DEC_WB/RegBank[27][3] ), 
        .B1(n17145), .B2(\pipeline/RegFile_DEC_WB/RegBank[26][3] ), .ZN(n16360) );
  AOI22_X1 U10702 ( .A1(n17146), .A2(\pipeline/RegFile_DEC_WB/RegBank[23][3] ), 
        .B1(n17147), .B2(\pipeline/RegFile_DEC_WB/RegBank[22][3] ), .ZN(n16361) );
  AOI22_X1 U10701 ( .A1(n17148), .A2(\pipeline/RegFile_DEC_WB/RegBank[21][3] ), 
        .B1(n17131), .B2(\pipeline/RegFile_DEC_WB/RegBank[20][3] ), .ZN(n16362) );
  AOI22_X1 U10700 ( .A1(n17128), .A2(\pipeline/RegFile_DEC_WB/RegBank[19][3] ), 
        .B1(n17134), .B2(\pipeline/RegFile_DEC_WB/RegBank[18][3] ), .ZN(n16363) );
  NAND4_X1 U10699 ( .A1(n16360), .A2(n16361), .A3(n16362), .A4(n16363), .ZN(
        n16349) );
  AOI22_X1 U10698 ( .A1(n17141), .A2(\pipeline/RegFile_DEC_WB/RegBank[17][3] ), 
        .B1(n17342), .B2(\pipeline/RegFile_DEC_WB/RegBank[16][3] ), .ZN(n16356) );
  AOI22_X1 U10697 ( .A1(n15916), .A2(\pipeline/RegFile_DEC_WB/RegBank[9][3] ), 
        .B1(n17139), .B2(\pipeline/RegFile_DEC_WB/RegBank[2][3] ), .ZN(n16357)
         );
  AOI22_X1 U10696 ( .A1(n17136), .A2(\pipeline/RegFile_DEC_WB/RegBank[12][3] ), 
        .B1(n15915), .B2(\pipeline/RegFile_DEC_WB/RegBank[11][3] ), .ZN(n16358) );
  AOI22_X1 U10695 ( .A1(n17140), .A2(\pipeline/RegFile_DEC_WB/RegBank[14][3] ), 
        .B1(n15913), .B2(\pipeline/RegFile_DEC_WB/RegBank[15][3] ), .ZN(n16359) );
  NAND4_X1 U10694 ( .A1(n16356), .A2(n16357), .A3(n16358), .A4(n16359), .ZN(
        n16350) );
  AOI22_X1 U10693 ( .A1(n17133), .A2(\pipeline/RegFile_DEC_WB/RegBank[13][3] ), 
        .B1(n15907), .B2(\pipeline/RegFile_DEC_WB/RegBank[4][3] ), .ZN(n16352)
         );
  AOI22_X1 U10692 ( .A1(n17335), .A2(\pipeline/RegFile_DEC_WB/RegBank[10][3] ), 
        .B1(n17144), .B2(\pipeline/RegFile_DEC_WB/RegBank[3][3] ), .ZN(n16353)
         );
  AOI22_X1 U10691 ( .A1(n17339), .A2(\pipeline/RegFile_DEC_WB/RegBank[6][3] ), 
        .B1(n17142), .B2(\pipeline/RegFile_DEC_WB/RegBank[7][3] ), .ZN(n16354)
         );
  AOI22_X1 U10690 ( .A1(n17337), .A2(\pipeline/RegFile_DEC_WB/RegBank[5][3] ), 
        .B1(n15901), .B2(\pipeline/RegFile_DEC_WB/RegBank[1][3] ), .ZN(n16355)
         );
  NAND4_X1 U10689 ( .A1(n16352), .A2(n16353), .A3(n16354), .A4(n16355), .ZN(
        n16351) );
  NOR4_X1 U10688 ( .A1(n16348), .A2(n16349), .A3(n16350), .A4(n16351), .ZN(
        n14939) );
  AOI22_X1 U10687 ( .A1(n17137), .A2(\pipeline/RegFile_DEC_WB/RegBank[31][2] ), 
        .B1(n17138), .B2(\pipeline/RegFile_DEC_WB/RegBank[30][2] ), .ZN(n16345) );
  AOI22_X1 U10686 ( .A1(n17130), .A2(\pipeline/RegFile_DEC_WB/RegBank[29][2] ), 
        .B1(n17129), .B2(\pipeline/RegFile_DEC_WB/RegBank[28][2] ), .ZN(n16346) );
  AOI222_X1 U10685 ( .A1(n17135), .A2(\pipeline/RegFile_DEC_WB/RegBank[8][2] ), 
        .B1(n17132), .B2(\pipeline/RegFile_DEC_WB/RegBank[25][2] ), .C1(n17127), .C2(\pipeline/RegFile_DEC_WB/RegBank[24][2] ), .ZN(n16347) );
  AOI22_X1 U10684 ( .A1(n17143), .A2(\pipeline/RegFile_DEC_WB/RegBank[27][2] ), 
        .B1(n17145), .B2(\pipeline/RegFile_DEC_WB/RegBank[26][2] ), .ZN(n16341) );
  AOI22_X1 U10683 ( .A1(n17146), .A2(\pipeline/RegFile_DEC_WB/RegBank[23][2] ), 
        .B1(n17147), .B2(\pipeline/RegFile_DEC_WB/RegBank[22][2] ), .ZN(n16342) );
  AOI22_X1 U10682 ( .A1(n17148), .A2(\pipeline/RegFile_DEC_WB/RegBank[21][2] ), 
        .B1(n17131), .B2(\pipeline/RegFile_DEC_WB/RegBank[20][2] ), .ZN(n16343) );
  AOI22_X1 U10681 ( .A1(n17128), .A2(\pipeline/RegFile_DEC_WB/RegBank[19][2] ), 
        .B1(n17134), .B2(\pipeline/RegFile_DEC_WB/RegBank[18][2] ), .ZN(n16344) );
  NAND4_X1 U10680 ( .A1(n16341), .A2(n16342), .A3(n16343), .A4(n16344), .ZN(
        n16330) );
  NOR2_X1 U10888 ( .A1(n16527), .A2(n16539), .ZN(n15919) );
  AOI22_X1 U10679 ( .A1(n17141), .A2(\pipeline/RegFile_DEC_WB/RegBank[17][2] ), 
        .B1(n15919), .B2(\pipeline/RegFile_DEC_WB/RegBank[16][2] ), .ZN(n16337) );
  AOI22_X1 U10678 ( .A1(n15916), .A2(\pipeline/RegFile_DEC_WB/RegBank[9][2] ), 
        .B1(n17139), .B2(\pipeline/RegFile_DEC_WB/RegBank[2][2] ), .ZN(n16338)
         );
  AOI22_X1 U10677 ( .A1(n17136), .A2(\pipeline/RegFile_DEC_WB/RegBank[12][2] ), 
        .B1(n15915), .B2(\pipeline/RegFile_DEC_WB/RegBank[11][2] ), .ZN(n16339) );
  AOI22_X1 U10676 ( .A1(n17140), .A2(\pipeline/RegFile_DEC_WB/RegBank[14][2] ), 
        .B1(n15913), .B2(\pipeline/RegFile_DEC_WB/RegBank[15][2] ), .ZN(n16340) );
  NAND4_X1 U10675 ( .A1(n16337), .A2(n16338), .A3(n16339), .A4(n16340), .ZN(
        n16331) );
  AOI22_X1 U10674 ( .A1(n17133), .A2(\pipeline/RegFile_DEC_WB/RegBank[13][2] ), 
        .B1(n15907), .B2(\pipeline/RegFile_DEC_WB/RegBank[4][2] ), .ZN(n16333)
         );
  NOR2_X1 U10873 ( .A1(n16533), .A2(n16532), .ZN(n15904) );
  AOI22_X1 U10673 ( .A1(n15904), .A2(\pipeline/RegFile_DEC_WB/RegBank[10][2] ), 
        .B1(n17144), .B2(\pipeline/RegFile_DEC_WB/RegBank[3][2] ), .ZN(n16334)
         );
  NOR2_X1 U10870 ( .A1(n16530), .A2(n16531), .ZN(n15902) );
  AOI22_X1 U10672 ( .A1(n15902), .A2(\pipeline/RegFile_DEC_WB/RegBank[6][2] ), 
        .B1(n17142), .B2(\pipeline/RegFile_DEC_WB/RegBank[7][2] ), .ZN(n16335)
         );
  AOI22_X1 U10671 ( .A1(n17345), .A2(\pipeline/RegFile_DEC_WB/RegBank[5][2] ), 
        .B1(n15901), .B2(\pipeline/RegFile_DEC_WB/RegBank[1][2] ), .ZN(n16336)
         );
  NAND4_X1 U10670 ( .A1(n16333), .A2(n16334), .A3(n16335), .A4(n16336), .ZN(
        n16332) );
  NOR4_X1 U10669 ( .A1(n16329), .A2(n16330), .A3(n16331), .A4(n16332), .ZN(
        n14941) );
  AOI22_X1 U10668 ( .A1(n17137), .A2(\pipeline/RegFile_DEC_WB/RegBank[31][1] ), 
        .B1(n17138), .B2(\pipeline/RegFile_DEC_WB/RegBank[30][1] ), .ZN(n16326) );
  AOI22_X1 U10667 ( .A1(n17130), .A2(\pipeline/RegFile_DEC_WB/RegBank[29][1] ), 
        .B1(n17129), .B2(\pipeline/RegFile_DEC_WB/RegBank[28][1] ), .ZN(n16327) );
  AOI222_X1 U10666 ( .A1(n17135), .A2(\pipeline/RegFile_DEC_WB/RegBank[8][1] ), 
        .B1(n17132), .B2(\pipeline/RegFile_DEC_WB/RegBank[25][1] ), .C1(n17127), .C2(\pipeline/RegFile_DEC_WB/RegBank[24][1] ), .ZN(n16328) );
  AOI22_X1 U10665 ( .A1(n17143), .A2(\pipeline/RegFile_DEC_WB/RegBank[27][1] ), 
        .B1(n17145), .B2(\pipeline/RegFile_DEC_WB/RegBank[26][1] ), .ZN(n16322) );
  AOI22_X1 U10664 ( .A1(n17146), .A2(\pipeline/RegFile_DEC_WB/RegBank[23][1] ), 
        .B1(n17147), .B2(\pipeline/RegFile_DEC_WB/RegBank[22][1] ), .ZN(n16323) );
  AOI22_X1 U10663 ( .A1(n17148), .A2(\pipeline/RegFile_DEC_WB/RegBank[21][1] ), 
        .B1(n17131), .B2(\pipeline/RegFile_DEC_WB/RegBank[20][1] ), .ZN(n16324) );
  AOI22_X1 U10662 ( .A1(n17128), .A2(\pipeline/RegFile_DEC_WB/RegBank[19][1] ), 
        .B1(n17134), .B2(\pipeline/RegFile_DEC_WB/RegBank[18][1] ), .ZN(n16325) );
  NAND4_X1 U10661 ( .A1(n16322), .A2(n16323), .A3(n16324), .A4(n16325), .ZN(
        n16311) );
  AOI22_X1 U10660 ( .A1(n17141), .A2(\pipeline/RegFile_DEC_WB/RegBank[17][1] ), 
        .B1(n15919), .B2(\pipeline/RegFile_DEC_WB/RegBank[16][1] ), .ZN(n16318) );
  AOI22_X1 U10659 ( .A1(n15916), .A2(\pipeline/RegFile_DEC_WB/RegBank[9][1] ), 
        .B1(n17139), .B2(\pipeline/RegFile_DEC_WB/RegBank[2][1] ), .ZN(n16319)
         );
  AOI22_X1 U10658 ( .A1(n17136), .A2(\pipeline/RegFile_DEC_WB/RegBank[12][1] ), 
        .B1(n15915), .B2(\pipeline/RegFile_DEC_WB/RegBank[11][1] ), .ZN(n16320) );
  AOI22_X1 U10657 ( .A1(n17140), .A2(\pipeline/RegFile_DEC_WB/RegBank[14][1] ), 
        .B1(n15913), .B2(\pipeline/RegFile_DEC_WB/RegBank[15][1] ), .ZN(n16321) );
  NAND4_X1 U10656 ( .A1(n16318), .A2(n16319), .A3(n16320), .A4(n16321), .ZN(
        n16312) );
  AOI22_X1 U10655 ( .A1(n17133), .A2(\pipeline/RegFile_DEC_WB/RegBank[13][1] ), 
        .B1(n15907), .B2(\pipeline/RegFile_DEC_WB/RegBank[4][1] ), .ZN(n16314)
         );
  AOI22_X1 U10654 ( .A1(n15904), .A2(\pipeline/RegFile_DEC_WB/RegBank[10][1] ), 
        .B1(n17144), .B2(\pipeline/RegFile_DEC_WB/RegBank[3][1] ), .ZN(n16315)
         );
  AOI22_X1 U10653 ( .A1(n15902), .A2(\pipeline/RegFile_DEC_WB/RegBank[6][1] ), 
        .B1(n17142), .B2(\pipeline/RegFile_DEC_WB/RegBank[7][1] ), .ZN(n16316)
         );
  AOI22_X1 U10652 ( .A1(n17345), .A2(\pipeline/RegFile_DEC_WB/RegBank[5][1] ), 
        .B1(n15901), .B2(\pipeline/RegFile_DEC_WB/RegBank[1][1] ), .ZN(n16317)
         );
  NAND4_X1 U10651 ( .A1(n16314), .A2(n16315), .A3(n16316), .A4(n16317), .ZN(
        n16313) );
  NOR4_X1 U10650 ( .A1(n16310), .A2(n16311), .A3(n16312), .A4(n16313), .ZN(
        n14943) );
  NAND4_X1 U10649 ( .A1(n14937), .A2(n14939), .A3(n14941), .A4(n14943), .ZN(
        n16309) );
  NOR4_X1 U10648 ( .A1(n15832), .A2(n15772), .A3(n15688), .A4(n16309), .ZN(
        n15999) );
  AOI22_X1 U10647 ( .A1(n17137), .A2(\pipeline/RegFile_DEC_WB/RegBank[31][18] ), .B1(n17138), .B2(\pipeline/RegFile_DEC_WB/RegBank[30][18] ), .ZN(n16306) );
  AOI22_X1 U10646 ( .A1(n17130), .A2(\pipeline/RegFile_DEC_WB/RegBank[29][18] ), .B1(n17129), .B2(\pipeline/RegFile_DEC_WB/RegBank[28][18] ), .ZN(n16307) );
  AOI222_X1 U10645 ( .A1(n17135), .A2(\pipeline/RegFile_DEC_WB/RegBank[8][18] ), .B1(n17132), .B2(\pipeline/RegFile_DEC_WB/RegBank[25][18] ), .C1(n17127), 
        .C2(\pipeline/RegFile_DEC_WB/RegBank[24][18] ), .ZN(n16308) );
  AOI22_X1 U10644 ( .A1(n17143), .A2(\pipeline/RegFile_DEC_WB/RegBank[27][18] ), .B1(n17145), .B2(\pipeline/RegFile_DEC_WB/RegBank[26][18] ), .ZN(n16302) );
  AOI22_X1 U10643 ( .A1(n17146), .A2(\pipeline/RegFile_DEC_WB/RegBank[23][18] ), .B1(n17147), .B2(\pipeline/RegFile_DEC_WB/RegBank[22][18] ), .ZN(n16303) );
  AOI22_X1 U10642 ( .A1(n17148), .A2(\pipeline/RegFile_DEC_WB/RegBank[21][18] ), .B1(n17131), .B2(\pipeline/RegFile_DEC_WB/RegBank[20][18] ), .ZN(n16304) );
  AOI22_X1 U10641 ( .A1(n17128), .A2(\pipeline/RegFile_DEC_WB/RegBank[19][18] ), .B1(n17134), .B2(\pipeline/RegFile_DEC_WB/RegBank[18][18] ), .ZN(n16305) );
  NAND4_X1 U10640 ( .A1(n16302), .A2(n16303), .A3(n16304), .A4(n16305), .ZN(
        n16291) );
  AOI22_X1 U10639 ( .A1(n17141), .A2(\pipeline/RegFile_DEC_WB/RegBank[17][18] ), .B1(n15919), .B2(\pipeline/RegFile_DEC_WB/RegBank[16][18] ), .ZN(n16298) );
  AOI22_X1 U10638 ( .A1(n15916), .A2(\pipeline/RegFile_DEC_WB/RegBank[9][18] ), 
        .B1(n17139), .B2(\pipeline/RegFile_DEC_WB/RegBank[2][18] ), .ZN(n16299) );
  AOI22_X1 U10637 ( .A1(n17136), .A2(\pipeline/RegFile_DEC_WB/RegBank[12][18] ), .B1(n15915), .B2(\pipeline/RegFile_DEC_WB/RegBank[11][18] ), .ZN(n16300) );
  AOI22_X1 U10636 ( .A1(n17140), .A2(\pipeline/RegFile_DEC_WB/RegBank[14][18] ), .B1(n15913), .B2(\pipeline/RegFile_DEC_WB/RegBank[15][18] ), .ZN(n16301) );
  NAND4_X1 U10635 ( .A1(n16298), .A2(n16299), .A3(n16300), .A4(n16301), .ZN(
        n16292) );
  AOI22_X1 U10634 ( .A1(n17133), .A2(\pipeline/RegFile_DEC_WB/RegBank[13][18] ), .B1(n15907), .B2(\pipeline/RegFile_DEC_WB/RegBank[4][18] ), .ZN(n16294) );
  AOI22_X1 U10633 ( .A1(n15904), .A2(\pipeline/RegFile_DEC_WB/RegBank[10][18] ), .B1(n17144), .B2(\pipeline/RegFile_DEC_WB/RegBank[3][18] ), .ZN(n16295) );
  AOI22_X1 U10632 ( .A1(n15902), .A2(\pipeline/RegFile_DEC_WB/RegBank[6][18] ), 
        .B1(n17142), .B2(\pipeline/RegFile_DEC_WB/RegBank[7][18] ), .ZN(n16296) );
  AOI22_X1 U10631 ( .A1(n17345), .A2(\pipeline/RegFile_DEC_WB/RegBank[5][18] ), 
        .B1(n15901), .B2(\pipeline/RegFile_DEC_WB/RegBank[1][18] ), .ZN(n16297) );
  NAND4_X1 U10630 ( .A1(n16294), .A2(n16295), .A3(n16296), .A4(n16297), .ZN(
        n16293) );
  NOR4_X1 U10629 ( .A1(n16290), .A2(n16291), .A3(n16292), .A4(n16293), .ZN(
        n14909) );
  AOI22_X1 U10628 ( .A1(n17137), .A2(\pipeline/RegFile_DEC_WB/RegBank[31][17] ), .B1(n17138), .B2(\pipeline/RegFile_DEC_WB/RegBank[30][17] ), .ZN(n16287) );
  AOI22_X1 U10627 ( .A1(n17130), .A2(\pipeline/RegFile_DEC_WB/RegBank[29][17] ), .B1(n17129), .B2(\pipeline/RegFile_DEC_WB/RegBank[28][17] ), .ZN(n16288) );
  AOI222_X1 U10626 ( .A1(n17135), .A2(\pipeline/RegFile_DEC_WB/RegBank[8][17] ), .B1(n17132), .B2(\pipeline/RegFile_DEC_WB/RegBank[25][17] ), .C1(n17127), 
        .C2(\pipeline/RegFile_DEC_WB/RegBank[24][17] ), .ZN(n16289) );
  AOI22_X1 U10625 ( .A1(n17143), .A2(\pipeline/RegFile_DEC_WB/RegBank[27][17] ), .B1(n17145), .B2(\pipeline/RegFile_DEC_WB/RegBank[26][17] ), .ZN(n16283) );
  AOI22_X1 U10624 ( .A1(n17146), .A2(\pipeline/RegFile_DEC_WB/RegBank[23][17] ), .B1(n17147), .B2(\pipeline/RegFile_DEC_WB/RegBank[22][17] ), .ZN(n16284) );
  AOI22_X1 U10623 ( .A1(n17148), .A2(\pipeline/RegFile_DEC_WB/RegBank[21][17] ), .B1(n17131), .B2(\pipeline/RegFile_DEC_WB/RegBank[20][17] ), .ZN(n16285) );
  AOI22_X1 U10622 ( .A1(n17128), .A2(\pipeline/RegFile_DEC_WB/RegBank[19][17] ), .B1(n17134), .B2(\pipeline/RegFile_DEC_WB/RegBank[18][17] ), .ZN(n16286) );
  NAND4_X1 U10621 ( .A1(n16283), .A2(n16284), .A3(n16285), .A4(n16286), .ZN(
        n16272) );
  AOI22_X1 U10620 ( .A1(n17141), .A2(\pipeline/RegFile_DEC_WB/RegBank[17][17] ), .B1(n17341), .B2(\pipeline/RegFile_DEC_WB/RegBank[16][17] ), .ZN(n16279) );
  AOI22_X1 U10619 ( .A1(n17388), .A2(\pipeline/RegFile_DEC_WB/RegBank[9][17] ), 
        .B1(n17139), .B2(\pipeline/RegFile_DEC_WB/RegBank[2][17] ), .ZN(n16280) );
  AOI22_X1 U10618 ( .A1(n17136), .A2(\pipeline/RegFile_DEC_WB/RegBank[12][17] ), .B1(n17389), .B2(\pipeline/RegFile_DEC_WB/RegBank[11][17] ), .ZN(n16281) );
  AOI22_X1 U10617 ( .A1(n17140), .A2(\pipeline/RegFile_DEC_WB/RegBank[14][17] ), .B1(n17390), .B2(\pipeline/RegFile_DEC_WB/RegBank[15][17] ), .ZN(n16282) );
  NAND4_X1 U10616 ( .A1(n16279), .A2(n16280), .A3(n16281), .A4(n16282), .ZN(
        n16273) );
  AOI22_X1 U10615 ( .A1(n17133), .A2(\pipeline/RegFile_DEC_WB/RegBank[13][17] ), .B1(n17392), .B2(\pipeline/RegFile_DEC_WB/RegBank[4][17] ), .ZN(n16275) );
  AOI22_X1 U10614 ( .A1(n17334), .A2(\pipeline/RegFile_DEC_WB/RegBank[10][17] ), .B1(n17144), .B2(\pipeline/RegFile_DEC_WB/RegBank[3][17] ), .ZN(n16276) );
  AOI22_X1 U10613 ( .A1(n17338), .A2(\pipeline/RegFile_DEC_WB/RegBank[6][17] ), 
        .B1(n17142), .B2(\pipeline/RegFile_DEC_WB/RegBank[7][17] ), .ZN(n16277) );
  AOI22_X1 U10612 ( .A1(n17336), .A2(\pipeline/RegFile_DEC_WB/RegBank[5][17] ), 
        .B1(n17391), .B2(\pipeline/RegFile_DEC_WB/RegBank[1][17] ), .ZN(n16278) );
  NAND4_X1 U10611 ( .A1(n16275), .A2(n16276), .A3(n16277), .A4(n16278), .ZN(
        n16274) );
  NOR4_X1 U10610 ( .A1(n16271), .A2(n16272), .A3(n16273), .A4(n16274), .ZN(
        n14911) );
  AOI22_X1 U10609 ( .A1(n15940), .A2(\pipeline/RegFile_DEC_WB/RegBank[31][16] ), .B1(n15941), .B2(\pipeline/RegFile_DEC_WB/RegBank[30][16] ), .ZN(n16268) );
  AOI22_X1 U10608 ( .A1(n15938), .A2(\pipeline/RegFile_DEC_WB/RegBank[29][16] ), .B1(n15939), .B2(\pipeline/RegFile_DEC_WB/RegBank[28][16] ), .ZN(n16269) );
  AOI222_X1 U10607 ( .A1(n15935), .A2(\pipeline/RegFile_DEC_WB/RegBank[8][16] ), .B1(n15936), .B2(\pipeline/RegFile_DEC_WB/RegBank[25][16] ), .C1(n15937), 
        .C2(\pipeline/RegFile_DEC_WB/RegBank[24][16] ), .ZN(n16270) );
  AOI22_X1 U10606 ( .A1(n15930), .A2(\pipeline/RegFile_DEC_WB/RegBank[27][16] ), .B1(n15931), .B2(\pipeline/RegFile_DEC_WB/RegBank[26][16] ), .ZN(n16264) );
  AOI22_X1 U10605 ( .A1(n15928), .A2(\pipeline/RegFile_DEC_WB/RegBank[23][16] ), .B1(n15929), .B2(\pipeline/RegFile_DEC_WB/RegBank[22][16] ), .ZN(n16265) );
  AOI22_X1 U10604 ( .A1(n15926), .A2(\pipeline/RegFile_DEC_WB/RegBank[21][16] ), .B1(n15927), .B2(\pipeline/RegFile_DEC_WB/RegBank[20][16] ), .ZN(n16266) );
  AOI22_X1 U10603 ( .A1(n15924), .A2(\pipeline/RegFile_DEC_WB/RegBank[19][16] ), .B1(n15925), .B2(\pipeline/RegFile_DEC_WB/RegBank[18][16] ), .ZN(n16267) );
  NAND4_X1 U10602 ( .A1(n16264), .A2(n16265), .A3(n16266), .A4(n16267), .ZN(
        n16253) );
  AOI22_X1 U10601 ( .A1(n15918), .A2(\pipeline/RegFile_DEC_WB/RegBank[17][16] ), .B1(n17342), .B2(\pipeline/RegFile_DEC_WB/RegBank[16][16] ), .ZN(n16260) );
  AOI22_X1 U10600 ( .A1(n15916), .A2(\pipeline/RegFile_DEC_WB/RegBank[9][16] ), 
        .B1(n15917), .B2(\pipeline/RegFile_DEC_WB/RegBank[2][16] ), .ZN(n16261) );
  AOI22_X1 U10599 ( .A1(n15914), .A2(\pipeline/RegFile_DEC_WB/RegBank[12][16] ), .B1(n15915), .B2(\pipeline/RegFile_DEC_WB/RegBank[11][16] ), .ZN(n16262) );
  AOI22_X1 U10598 ( .A1(n15912), .A2(\pipeline/RegFile_DEC_WB/RegBank[14][16] ), .B1(n15913), .B2(\pipeline/RegFile_DEC_WB/RegBank[15][16] ), .ZN(n16263) );
  NAND4_X1 U10597 ( .A1(n16260), .A2(n16261), .A3(n16262), .A4(n16263), .ZN(
        n16254) );
  AOI22_X1 U10596 ( .A1(n15906), .A2(\pipeline/RegFile_DEC_WB/RegBank[13][16] ), .B1(n15907), .B2(\pipeline/RegFile_DEC_WB/RegBank[4][16] ), .ZN(n16256) );
  AOI22_X1 U10595 ( .A1(n17335), .A2(\pipeline/RegFile_DEC_WB/RegBank[10][16] ), .B1(n15905), .B2(\pipeline/RegFile_DEC_WB/RegBank[3][16] ), .ZN(n16257) );
  AOI22_X1 U10594 ( .A1(n17339), .A2(\pipeline/RegFile_DEC_WB/RegBank[6][16] ), 
        .B1(n15903), .B2(\pipeline/RegFile_DEC_WB/RegBank[7][16] ), .ZN(n16258) );
  AOI22_X1 U10593 ( .A1(n17337), .A2(\pipeline/RegFile_DEC_WB/RegBank[5][16] ), 
        .B1(n15901), .B2(\pipeline/RegFile_DEC_WB/RegBank[1][16] ), .ZN(n16259) );
  NAND4_X1 U10592 ( .A1(n16256), .A2(n16257), .A3(n16258), .A4(n16259), .ZN(
        n16255) );
  NOR4_X1 U10591 ( .A1(n16252), .A2(n16253), .A3(n16254), .A4(n16255), .ZN(
        n14913) );
  AOI22_X1 U10590 ( .A1(n15940), .A2(\pipeline/RegFile_DEC_WB/RegBank[31][15] ), .B1(n15941), .B2(\pipeline/RegFile_DEC_WB/RegBank[30][15] ), .ZN(n16249) );
  AOI22_X1 U10589 ( .A1(n15938), .A2(\pipeline/RegFile_DEC_WB/RegBank[29][15] ), .B1(n15939), .B2(\pipeline/RegFile_DEC_WB/RegBank[28][15] ), .ZN(n16250) );
  AOI222_X1 U10588 ( .A1(n15935), .A2(\pipeline/RegFile_DEC_WB/RegBank[8][15] ), .B1(n15936), .B2(\pipeline/RegFile_DEC_WB/RegBank[25][15] ), .C1(n15937), 
        .C2(\pipeline/RegFile_DEC_WB/RegBank[24][15] ), .ZN(n16251) );
  AOI22_X1 U10587 ( .A1(n15930), .A2(\pipeline/RegFile_DEC_WB/RegBank[27][15] ), .B1(n15931), .B2(\pipeline/RegFile_DEC_WB/RegBank[26][15] ), .ZN(n16245) );
  AOI22_X1 U10586 ( .A1(n15928), .A2(\pipeline/RegFile_DEC_WB/RegBank[23][15] ), .B1(n15929), .B2(\pipeline/RegFile_DEC_WB/RegBank[22][15] ), .ZN(n16246) );
  AOI22_X1 U10585 ( .A1(n15926), .A2(\pipeline/RegFile_DEC_WB/RegBank[21][15] ), .B1(n15927), .B2(\pipeline/RegFile_DEC_WB/RegBank[20][15] ), .ZN(n16247) );
  AOI22_X1 U10584 ( .A1(n15924), .A2(\pipeline/RegFile_DEC_WB/RegBank[19][15] ), .B1(n15925), .B2(\pipeline/RegFile_DEC_WB/RegBank[18][15] ), .ZN(n16248) );
  NAND4_X1 U10583 ( .A1(n16245), .A2(n16246), .A3(n16247), .A4(n16248), .ZN(
        n16234) );
  AOI22_X1 U10582 ( .A1(n15918), .A2(\pipeline/RegFile_DEC_WB/RegBank[17][15] ), .B1(n17342), .B2(\pipeline/RegFile_DEC_WB/RegBank[16][15] ), .ZN(n16241) );
  AOI22_X1 U10581 ( .A1(n15916), .A2(\pipeline/RegFile_DEC_WB/RegBank[9][15] ), 
        .B1(n15917), .B2(\pipeline/RegFile_DEC_WB/RegBank[2][15] ), .ZN(n16242) );
  AOI22_X1 U10580 ( .A1(n15914), .A2(\pipeline/RegFile_DEC_WB/RegBank[12][15] ), .B1(n15915), .B2(\pipeline/RegFile_DEC_WB/RegBank[11][15] ), .ZN(n16243) );
  AOI22_X1 U10579 ( .A1(n15912), .A2(\pipeline/RegFile_DEC_WB/RegBank[14][15] ), .B1(n15913), .B2(\pipeline/RegFile_DEC_WB/RegBank[15][15] ), .ZN(n16244) );
  NAND4_X1 U10578 ( .A1(n16241), .A2(n16242), .A3(n16243), .A4(n16244), .ZN(
        n16235) );
  AOI22_X1 U10577 ( .A1(n15906), .A2(\pipeline/RegFile_DEC_WB/RegBank[13][15] ), .B1(n15907), .B2(\pipeline/RegFile_DEC_WB/RegBank[4][15] ), .ZN(n16237) );
  AOI22_X1 U10576 ( .A1(n17335), .A2(\pipeline/RegFile_DEC_WB/RegBank[10][15] ), .B1(n15905), .B2(\pipeline/RegFile_DEC_WB/RegBank[3][15] ), .ZN(n16238) );
  AOI22_X1 U10575 ( .A1(n17339), .A2(\pipeline/RegFile_DEC_WB/RegBank[6][15] ), 
        .B1(n15903), .B2(\pipeline/RegFile_DEC_WB/RegBank[7][15] ), .ZN(n16239) );
  AOI22_X1 U10574 ( .A1(n17337), .A2(\pipeline/RegFile_DEC_WB/RegBank[5][15] ), 
        .B1(n15901), .B2(\pipeline/RegFile_DEC_WB/RegBank[1][15] ), .ZN(n16240) );
  NAND4_X1 U10573 ( .A1(n16237), .A2(n16238), .A3(n16239), .A4(n16240), .ZN(
        n16236) );
  NOR4_X1 U10572 ( .A1(n16233), .A2(n16234), .A3(n16235), .A4(n16236), .ZN(
        n14915) );
  NAND4_X1 U10571 ( .A1(n14909), .A2(n14911), .A3(n14913), .A4(n14915), .ZN(
        n16001) );
  AOI22_X1 U10570 ( .A1(n17137), .A2(\pipeline/RegFile_DEC_WB/RegBank[31][22] ), .B1(n17138), .B2(\pipeline/RegFile_DEC_WB/RegBank[30][22] ), .ZN(n16230) );
  AOI22_X1 U10569 ( .A1(n17130), .A2(\pipeline/RegFile_DEC_WB/RegBank[29][22] ), .B1(n17129), .B2(\pipeline/RegFile_DEC_WB/RegBank[28][22] ), .ZN(n16231) );
  AOI222_X1 U10568 ( .A1(n17135), .A2(\pipeline/RegFile_DEC_WB/RegBank[8][22] ), .B1(n17132), .B2(\pipeline/RegFile_DEC_WB/RegBank[25][22] ), .C1(n17127), 
        .C2(\pipeline/RegFile_DEC_WB/RegBank[24][22] ), .ZN(n16232) );
  AOI22_X1 U10567 ( .A1(n17143), .A2(\pipeline/RegFile_DEC_WB/RegBank[27][22] ), .B1(n17145), .B2(\pipeline/RegFile_DEC_WB/RegBank[26][22] ), .ZN(n16226) );
  AOI22_X1 U10566 ( .A1(n17146), .A2(\pipeline/RegFile_DEC_WB/RegBank[23][22] ), .B1(n17147), .B2(\pipeline/RegFile_DEC_WB/RegBank[22][22] ), .ZN(n16227) );
  AOI22_X1 U10565 ( .A1(n17148), .A2(\pipeline/RegFile_DEC_WB/RegBank[21][22] ), .B1(n17131), .B2(\pipeline/RegFile_DEC_WB/RegBank[20][22] ), .ZN(n16228) );
  AOI22_X1 U10564 ( .A1(n17128), .A2(\pipeline/RegFile_DEC_WB/RegBank[19][22] ), .B1(n17134), .B2(\pipeline/RegFile_DEC_WB/RegBank[18][22] ), .ZN(n16229) );
  NAND4_X1 U10563 ( .A1(n16226), .A2(n16227), .A3(n16228), .A4(n16229), .ZN(
        n16215) );
  AOI22_X1 U10562 ( .A1(n17141), .A2(\pipeline/RegFile_DEC_WB/RegBank[17][22] ), .B1(n15919), .B2(\pipeline/RegFile_DEC_WB/RegBank[16][22] ), .ZN(n16222) );
  AOI22_X1 U10561 ( .A1(n15916), .A2(\pipeline/RegFile_DEC_WB/RegBank[9][22] ), 
        .B1(n17139), .B2(\pipeline/RegFile_DEC_WB/RegBank[2][22] ), .ZN(n16223) );
  AOI22_X1 U10560 ( .A1(n17136), .A2(\pipeline/RegFile_DEC_WB/RegBank[12][22] ), .B1(n15915), .B2(\pipeline/RegFile_DEC_WB/RegBank[11][22] ), .ZN(n16224) );
  AOI22_X1 U10559 ( .A1(n17140), .A2(\pipeline/RegFile_DEC_WB/RegBank[14][22] ), .B1(n15913), .B2(\pipeline/RegFile_DEC_WB/RegBank[15][22] ), .ZN(n16225) );
  NAND4_X1 U10558 ( .A1(n16222), .A2(n16223), .A3(n16224), .A4(n16225), .ZN(
        n16216) );
  AOI22_X1 U10557 ( .A1(n17133), .A2(\pipeline/RegFile_DEC_WB/RegBank[13][22] ), .B1(n15907), .B2(\pipeline/RegFile_DEC_WB/RegBank[4][22] ), .ZN(n16218) );
  AOI22_X1 U10556 ( .A1(n15904), .A2(\pipeline/RegFile_DEC_WB/RegBank[10][22] ), .B1(n17144), .B2(\pipeline/RegFile_DEC_WB/RegBank[3][22] ), .ZN(n16219) );
  AOI22_X1 U10555 ( .A1(n15902), .A2(\pipeline/RegFile_DEC_WB/RegBank[6][22] ), 
        .B1(n17142), .B2(\pipeline/RegFile_DEC_WB/RegBank[7][22] ), .ZN(n16220) );
  AOI22_X1 U10554 ( .A1(n17345), .A2(\pipeline/RegFile_DEC_WB/RegBank[5][22] ), 
        .B1(n15901), .B2(\pipeline/RegFile_DEC_WB/RegBank[1][22] ), .ZN(n16221) );
  NAND4_X1 U10553 ( .A1(n16218), .A2(n16219), .A3(n16220), .A4(n16221), .ZN(
        n16217) );
  NOR4_X1 U10552 ( .A1(n16214), .A2(n16215), .A3(n16216), .A4(n16217), .ZN(
        n14901) );
  AOI22_X1 U10551 ( .A1(n17137), .A2(\pipeline/RegFile_DEC_WB/RegBank[31][21] ), .B1(n17138), .B2(\pipeline/RegFile_DEC_WB/RegBank[30][21] ), .ZN(n16211) );
  AOI22_X1 U10550 ( .A1(n17130), .A2(\pipeline/RegFile_DEC_WB/RegBank[29][21] ), .B1(n17129), .B2(\pipeline/RegFile_DEC_WB/RegBank[28][21] ), .ZN(n16212) );
  AOI222_X1 U10549 ( .A1(n17135), .A2(\pipeline/RegFile_DEC_WB/RegBank[8][21] ), .B1(n17132), .B2(\pipeline/RegFile_DEC_WB/RegBank[25][21] ), .C1(n17127), 
        .C2(\pipeline/RegFile_DEC_WB/RegBank[24][21] ), .ZN(n16213) );
  AOI22_X1 U10548 ( .A1(n17143), .A2(\pipeline/RegFile_DEC_WB/RegBank[27][21] ), .B1(n17145), .B2(\pipeline/RegFile_DEC_WB/RegBank[26][21] ), .ZN(n16207) );
  AOI22_X1 U10547 ( .A1(n17146), .A2(\pipeline/RegFile_DEC_WB/RegBank[23][21] ), .B1(n17147), .B2(\pipeline/RegFile_DEC_WB/RegBank[22][21] ), .ZN(n16208) );
  AOI22_X1 U10546 ( .A1(n17148), .A2(\pipeline/RegFile_DEC_WB/RegBank[21][21] ), .B1(n17131), .B2(\pipeline/RegFile_DEC_WB/RegBank[20][21] ), .ZN(n16209) );
  AOI22_X1 U10545 ( .A1(n17128), .A2(\pipeline/RegFile_DEC_WB/RegBank[19][21] ), .B1(n17134), .B2(\pipeline/RegFile_DEC_WB/RegBank[18][21] ), .ZN(n16210) );
  NAND4_X1 U10544 ( .A1(n16207), .A2(n16208), .A3(n16209), .A4(n16210), .ZN(
        n16196) );
  AOI22_X1 U10543 ( .A1(n17141), .A2(\pipeline/RegFile_DEC_WB/RegBank[17][21] ), .B1(n15919), .B2(\pipeline/RegFile_DEC_WB/RegBank[16][21] ), .ZN(n16203) );
  AOI22_X1 U10542 ( .A1(n15916), .A2(\pipeline/RegFile_DEC_WB/RegBank[9][21] ), 
        .B1(n17139), .B2(\pipeline/RegFile_DEC_WB/RegBank[2][21] ), .ZN(n16204) );
  AOI22_X1 U10541 ( .A1(n17136), .A2(\pipeline/RegFile_DEC_WB/RegBank[12][21] ), .B1(n15915), .B2(\pipeline/RegFile_DEC_WB/RegBank[11][21] ), .ZN(n16205) );
  AOI22_X1 U10540 ( .A1(n17140), .A2(\pipeline/RegFile_DEC_WB/RegBank[14][21] ), .B1(n15913), .B2(\pipeline/RegFile_DEC_WB/RegBank[15][21] ), .ZN(n16206) );
  NAND4_X1 U10539 ( .A1(n16203), .A2(n16204), .A3(n16205), .A4(n16206), .ZN(
        n16197) );
  AOI22_X1 U10538 ( .A1(n17133), .A2(\pipeline/RegFile_DEC_WB/RegBank[13][21] ), .B1(n15907), .B2(\pipeline/RegFile_DEC_WB/RegBank[4][21] ), .ZN(n16199) );
  AOI22_X1 U10537 ( .A1(n15904), .A2(\pipeline/RegFile_DEC_WB/RegBank[10][21] ), .B1(n17144), .B2(\pipeline/RegFile_DEC_WB/RegBank[3][21] ), .ZN(n16200) );
  AOI22_X1 U10536 ( .A1(n15902), .A2(\pipeline/RegFile_DEC_WB/RegBank[6][21] ), 
        .B1(n17142), .B2(\pipeline/RegFile_DEC_WB/RegBank[7][21] ), .ZN(n16201) );
  AOI22_X1 U10535 ( .A1(n17345), .A2(\pipeline/RegFile_DEC_WB/RegBank[5][21] ), 
        .B1(n15901), .B2(\pipeline/RegFile_DEC_WB/RegBank[1][21] ), .ZN(n16202) );
  NAND4_X1 U10534 ( .A1(n16199), .A2(n16200), .A3(n16201), .A4(n16202), .ZN(
        n16198) );
  NOR4_X1 U10533 ( .A1(n16195), .A2(n16196), .A3(n16197), .A4(n16198), .ZN(
        n14903) );
  AOI22_X1 U10532 ( .A1(n17137), .A2(\pipeline/RegFile_DEC_WB/RegBank[31][20] ), .B1(n17138), .B2(\pipeline/RegFile_DEC_WB/RegBank[30][20] ), .ZN(n16192) );
  AOI22_X1 U10531 ( .A1(n17130), .A2(\pipeline/RegFile_DEC_WB/RegBank[29][20] ), .B1(n17129), .B2(\pipeline/RegFile_DEC_WB/RegBank[28][20] ), .ZN(n16193) );
  AOI222_X1 U10530 ( .A1(n17135), .A2(\pipeline/RegFile_DEC_WB/RegBank[8][20] ), .B1(n17132), .B2(\pipeline/RegFile_DEC_WB/RegBank[25][20] ), .C1(n17127), 
        .C2(\pipeline/RegFile_DEC_WB/RegBank[24][20] ), .ZN(n16194) );
  AOI22_X1 U10529 ( .A1(n17143), .A2(\pipeline/RegFile_DEC_WB/RegBank[27][20] ), .B1(n17145), .B2(\pipeline/RegFile_DEC_WB/RegBank[26][20] ), .ZN(n16188) );
  AOI22_X1 U10528 ( .A1(n17146), .A2(\pipeline/RegFile_DEC_WB/RegBank[23][20] ), .B1(n17147), .B2(\pipeline/RegFile_DEC_WB/RegBank[22][20] ), .ZN(n16189) );
  AOI22_X1 U10527 ( .A1(n17148), .A2(\pipeline/RegFile_DEC_WB/RegBank[21][20] ), .B1(n17131), .B2(\pipeline/RegFile_DEC_WB/RegBank[20][20] ), .ZN(n16190) );
  AOI22_X1 U10526 ( .A1(n17128), .A2(\pipeline/RegFile_DEC_WB/RegBank[19][20] ), .B1(n17134), .B2(\pipeline/RegFile_DEC_WB/RegBank[18][20] ), .ZN(n16191) );
  NAND4_X1 U10525 ( .A1(n16188), .A2(n16189), .A3(n16190), .A4(n16191), .ZN(
        n16177) );
  AOI22_X1 U10524 ( .A1(n17141), .A2(\pipeline/RegFile_DEC_WB/RegBank[17][20] ), .B1(n15919), .B2(\pipeline/RegFile_DEC_WB/RegBank[16][20] ), .ZN(n16184) );
  AOI22_X1 U10523 ( .A1(n15916), .A2(\pipeline/RegFile_DEC_WB/RegBank[9][20] ), 
        .B1(n17139), .B2(\pipeline/RegFile_DEC_WB/RegBank[2][20] ), .ZN(n16185) );
  AOI22_X1 U10522 ( .A1(n17136), .A2(\pipeline/RegFile_DEC_WB/RegBank[12][20] ), .B1(n15915), .B2(\pipeline/RegFile_DEC_WB/RegBank[11][20] ), .ZN(n16186) );
  AOI22_X1 U10521 ( .A1(n17140), .A2(\pipeline/RegFile_DEC_WB/RegBank[14][20] ), .B1(n15913), .B2(\pipeline/RegFile_DEC_WB/RegBank[15][20] ), .ZN(n16187) );
  NAND4_X1 U10520 ( .A1(n16184), .A2(n16185), .A3(n16186), .A4(n16187), .ZN(
        n16178) );
  AOI22_X1 U10519 ( .A1(n17133), .A2(\pipeline/RegFile_DEC_WB/RegBank[13][20] ), .B1(n15907), .B2(\pipeline/RegFile_DEC_WB/RegBank[4][20] ), .ZN(n16180) );
  AOI22_X1 U10518 ( .A1(n15904), .A2(\pipeline/RegFile_DEC_WB/RegBank[10][20] ), .B1(n17144), .B2(\pipeline/RegFile_DEC_WB/RegBank[3][20] ), .ZN(n16181) );
  AOI22_X1 U10517 ( .A1(n15902), .A2(\pipeline/RegFile_DEC_WB/RegBank[6][20] ), 
        .B1(n17142), .B2(\pipeline/RegFile_DEC_WB/RegBank[7][20] ), .ZN(n16182) );
  AOI22_X1 U10516 ( .A1(n17345), .A2(\pipeline/RegFile_DEC_WB/RegBank[5][20] ), 
        .B1(n15901), .B2(\pipeline/RegFile_DEC_WB/RegBank[1][20] ), .ZN(n16183) );
  NAND4_X1 U10515 ( .A1(n16180), .A2(n16181), .A3(n16182), .A4(n16183), .ZN(
        n16179) );
  NOR4_X1 U10514 ( .A1(n16176), .A2(n16177), .A3(n16178), .A4(n16179), .ZN(
        n14905) );
  AOI22_X1 U10513 ( .A1(n15940), .A2(\pipeline/RegFile_DEC_WB/RegBank[31][19] ), .B1(n15941), .B2(\pipeline/RegFile_DEC_WB/RegBank[30][19] ), .ZN(n16173) );
  AOI22_X1 U10512 ( .A1(n15938), .A2(\pipeline/RegFile_DEC_WB/RegBank[29][19] ), .B1(n15939), .B2(\pipeline/RegFile_DEC_WB/RegBank[28][19] ), .ZN(n16174) );
  AOI222_X1 U10511 ( .A1(n15935), .A2(\pipeline/RegFile_DEC_WB/RegBank[8][19] ), .B1(n15936), .B2(\pipeline/RegFile_DEC_WB/RegBank[25][19] ), .C1(n15937), 
        .C2(\pipeline/RegFile_DEC_WB/RegBank[24][19] ), .ZN(n16175) );
  AOI22_X1 U10510 ( .A1(n15930), .A2(\pipeline/RegFile_DEC_WB/RegBank[27][19] ), .B1(n15931), .B2(\pipeline/RegFile_DEC_WB/RegBank[26][19] ), .ZN(n16169) );
  AOI22_X1 U10509 ( .A1(n15928), .A2(\pipeline/RegFile_DEC_WB/RegBank[23][19] ), .B1(n15929), .B2(\pipeline/RegFile_DEC_WB/RegBank[22][19] ), .ZN(n16170) );
  AOI22_X1 U10508 ( .A1(n15926), .A2(\pipeline/RegFile_DEC_WB/RegBank[21][19] ), .B1(n15927), .B2(\pipeline/RegFile_DEC_WB/RegBank[20][19] ), .ZN(n16171) );
  AOI22_X1 U10507 ( .A1(n15924), .A2(\pipeline/RegFile_DEC_WB/RegBank[19][19] ), .B1(n15925), .B2(\pipeline/RegFile_DEC_WB/RegBank[18][19] ), .ZN(n16172) );
  NAND4_X1 U10506 ( .A1(n16169), .A2(n16170), .A3(n16171), .A4(n16172), .ZN(
        n16158) );
  AOI22_X1 U10505 ( .A1(n15918), .A2(\pipeline/RegFile_DEC_WB/RegBank[17][19] ), .B1(n15919), .B2(\pipeline/RegFile_DEC_WB/RegBank[16][19] ), .ZN(n16165) );
  AOI22_X1 U10504 ( .A1(n15916), .A2(\pipeline/RegFile_DEC_WB/RegBank[9][19] ), 
        .B1(n15917), .B2(\pipeline/RegFile_DEC_WB/RegBank[2][19] ), .ZN(n16166) );
  AOI22_X1 U10503 ( .A1(n15914), .A2(\pipeline/RegFile_DEC_WB/RegBank[12][19] ), .B1(n15915), .B2(\pipeline/RegFile_DEC_WB/RegBank[11][19] ), .ZN(n16167) );
  AOI22_X1 U10502 ( .A1(n15912), .A2(\pipeline/RegFile_DEC_WB/RegBank[14][19] ), .B1(n15913), .B2(\pipeline/RegFile_DEC_WB/RegBank[15][19] ), .ZN(n16168) );
  NAND4_X1 U10501 ( .A1(n16165), .A2(n16166), .A3(n16167), .A4(n16168), .ZN(
        n16159) );
  AOI22_X1 U10500 ( .A1(n15906), .A2(\pipeline/RegFile_DEC_WB/RegBank[13][19] ), .B1(n15907), .B2(\pipeline/RegFile_DEC_WB/RegBank[4][19] ), .ZN(n16161) );
  AOI22_X1 U10499 ( .A1(n15904), .A2(\pipeline/RegFile_DEC_WB/RegBank[10][19] ), .B1(n15905), .B2(\pipeline/RegFile_DEC_WB/RegBank[3][19] ), .ZN(n16162) );
  AOI22_X1 U10498 ( .A1(n15902), .A2(\pipeline/RegFile_DEC_WB/RegBank[6][19] ), 
        .B1(n15903), .B2(\pipeline/RegFile_DEC_WB/RegBank[7][19] ), .ZN(n16163) );
  AOI22_X1 U10497 ( .A1(n17345), .A2(\pipeline/RegFile_DEC_WB/RegBank[5][19] ), 
        .B1(n15901), .B2(\pipeline/RegFile_DEC_WB/RegBank[1][19] ), .ZN(n16164) );
  NAND4_X1 U10496 ( .A1(n16161), .A2(n16162), .A3(n16163), .A4(n16164), .ZN(
        n16160) );
  NOR4_X1 U10495 ( .A1(n16157), .A2(n16158), .A3(n16159), .A4(n16160), .ZN(
        n14907) );
  NAND4_X1 U10494 ( .A1(n14901), .A2(n14903), .A3(n14905), .A4(n14907), .ZN(
        n16002) );
  AOI22_X1 U10493 ( .A1(n17137), .A2(\pipeline/RegFile_DEC_WB/RegBank[31][10] ), .B1(n17138), .B2(\pipeline/RegFile_DEC_WB/RegBank[30][10] ), .ZN(n16154) );
  AOI22_X1 U10492 ( .A1(n17130), .A2(\pipeline/RegFile_DEC_WB/RegBank[29][10] ), .B1(n17129), .B2(\pipeline/RegFile_DEC_WB/RegBank[28][10] ), .ZN(n16155) );
  AOI222_X1 U10491 ( .A1(n17135), .A2(\pipeline/RegFile_DEC_WB/RegBank[8][10] ), .B1(n17132), .B2(\pipeline/RegFile_DEC_WB/RegBank[25][10] ), .C1(n17127), 
        .C2(\pipeline/RegFile_DEC_WB/RegBank[24][10] ), .ZN(n16156) );
  AOI22_X1 U10490 ( .A1(n17143), .A2(\pipeline/RegFile_DEC_WB/RegBank[27][10] ), .B1(n17145), .B2(\pipeline/RegFile_DEC_WB/RegBank[26][10] ), .ZN(n16150) );
  AOI22_X1 U10489 ( .A1(n17146), .A2(\pipeline/RegFile_DEC_WB/RegBank[23][10] ), .B1(n17147), .B2(\pipeline/RegFile_DEC_WB/RegBank[22][10] ), .ZN(n16151) );
  AOI22_X1 U10488 ( .A1(n17148), .A2(\pipeline/RegFile_DEC_WB/RegBank[21][10] ), .B1(n17131), .B2(\pipeline/RegFile_DEC_WB/RegBank[20][10] ), .ZN(n16152) );
  AOI22_X1 U10487 ( .A1(n17128), .A2(\pipeline/RegFile_DEC_WB/RegBank[19][10] ), .B1(n17134), .B2(\pipeline/RegFile_DEC_WB/RegBank[18][10] ), .ZN(n16153) );
  NAND4_X1 U10486 ( .A1(n16150), .A2(n16151), .A3(n16152), .A4(n16153), .ZN(
        n16139) );
  AOI22_X1 U10485 ( .A1(n17141), .A2(\pipeline/RegFile_DEC_WB/RegBank[17][10] ), .B1(n15919), .B2(\pipeline/RegFile_DEC_WB/RegBank[16][10] ), .ZN(n16146) );
  AOI22_X1 U10484 ( .A1(n15916), .A2(\pipeline/RegFile_DEC_WB/RegBank[9][10] ), 
        .B1(n17139), .B2(\pipeline/RegFile_DEC_WB/RegBank[2][10] ), .ZN(n16147) );
  AOI22_X1 U10483 ( .A1(n17136), .A2(\pipeline/RegFile_DEC_WB/RegBank[12][10] ), .B1(n15915), .B2(\pipeline/RegFile_DEC_WB/RegBank[11][10] ), .ZN(n16148) );
  AOI22_X1 U10482 ( .A1(n17140), .A2(\pipeline/RegFile_DEC_WB/RegBank[14][10] ), .B1(n15913), .B2(\pipeline/RegFile_DEC_WB/RegBank[15][10] ), .ZN(n16149) );
  NAND4_X1 U10481 ( .A1(n16146), .A2(n16147), .A3(n16148), .A4(n16149), .ZN(
        n16140) );
  AOI22_X1 U10480 ( .A1(n17133), .A2(\pipeline/RegFile_DEC_WB/RegBank[13][10] ), .B1(n15907), .B2(\pipeline/RegFile_DEC_WB/RegBank[4][10] ), .ZN(n16142) );
  AOI22_X1 U10479 ( .A1(n15904), .A2(\pipeline/RegFile_DEC_WB/RegBank[10][10] ), .B1(n17144), .B2(\pipeline/RegFile_DEC_WB/RegBank[3][10] ), .ZN(n16143) );
  AOI22_X1 U10478 ( .A1(n15902), .A2(\pipeline/RegFile_DEC_WB/RegBank[6][10] ), 
        .B1(n17142), .B2(\pipeline/RegFile_DEC_WB/RegBank[7][10] ), .ZN(n16144) );
  AOI22_X1 U10477 ( .A1(n17345), .A2(\pipeline/RegFile_DEC_WB/RegBank[5][10] ), 
        .B1(n15901), .B2(\pipeline/RegFile_DEC_WB/RegBank[1][10] ), .ZN(n16145) );
  NAND4_X1 U10476 ( .A1(n16142), .A2(n16143), .A3(n16144), .A4(n16145), .ZN(
        n16141) );
  NOR4_X1 U10475 ( .A1(n16138), .A2(n16139), .A3(n16140), .A4(n16141), .ZN(
        n14925) );
  AOI22_X1 U10474 ( .A1(n17137), .A2(\pipeline/RegFile_DEC_WB/RegBank[31][9] ), 
        .B1(n17138), .B2(\pipeline/RegFile_DEC_WB/RegBank[30][9] ), .ZN(n16135) );
  AOI22_X1 U10473 ( .A1(n17130), .A2(\pipeline/RegFile_DEC_WB/RegBank[29][9] ), 
        .B1(n17129), .B2(\pipeline/RegFile_DEC_WB/RegBank[28][9] ), .ZN(n16136) );
  AOI222_X1 U10472 ( .A1(n17135), .A2(\pipeline/RegFile_DEC_WB/RegBank[8][9] ), 
        .B1(n17132), .B2(\pipeline/RegFile_DEC_WB/RegBank[25][9] ), .C1(n17127), .C2(\pipeline/RegFile_DEC_WB/RegBank[24][9] ), .ZN(n16137) );
  AOI22_X1 U10471 ( .A1(n17143), .A2(\pipeline/RegFile_DEC_WB/RegBank[27][9] ), 
        .B1(n17145), .B2(\pipeline/RegFile_DEC_WB/RegBank[26][9] ), .ZN(n16131) );
  AOI22_X1 U10470 ( .A1(n17146), .A2(\pipeline/RegFile_DEC_WB/RegBank[23][9] ), 
        .B1(n17147), .B2(\pipeline/RegFile_DEC_WB/RegBank[22][9] ), .ZN(n16132) );
  AOI22_X1 U10469 ( .A1(n17148), .A2(\pipeline/RegFile_DEC_WB/RegBank[21][9] ), 
        .B1(n17131), .B2(\pipeline/RegFile_DEC_WB/RegBank[20][9] ), .ZN(n16133) );
  AOI22_X1 U10468 ( .A1(n17128), .A2(\pipeline/RegFile_DEC_WB/RegBank[19][9] ), 
        .B1(n17134), .B2(\pipeline/RegFile_DEC_WB/RegBank[18][9] ), .ZN(n16134) );
  NAND4_X1 U10467 ( .A1(n16131), .A2(n16132), .A3(n16133), .A4(n16134), .ZN(
        n16120) );
  AOI22_X1 U10466 ( .A1(n17141), .A2(\pipeline/RegFile_DEC_WB/RegBank[17][9] ), 
        .B1(n17341), .B2(\pipeline/RegFile_DEC_WB/RegBank[16][9] ), .ZN(n16127) );
  AOI22_X1 U10465 ( .A1(n17388), .A2(\pipeline/RegFile_DEC_WB/RegBank[9][9] ), 
        .B1(n17139), .B2(\pipeline/RegFile_DEC_WB/RegBank[2][9] ), .ZN(n16128)
         );
  AOI22_X1 U10464 ( .A1(n17136), .A2(\pipeline/RegFile_DEC_WB/RegBank[12][9] ), 
        .B1(n17389), .B2(\pipeline/RegFile_DEC_WB/RegBank[11][9] ), .ZN(n16129) );
  AOI22_X1 U10463 ( .A1(n17140), .A2(\pipeline/RegFile_DEC_WB/RegBank[14][9] ), 
        .B1(n17390), .B2(\pipeline/RegFile_DEC_WB/RegBank[15][9] ), .ZN(n16130) );
  NAND4_X1 U10462 ( .A1(n16127), .A2(n16128), .A3(n16129), .A4(n16130), .ZN(
        n16121) );
  AOI22_X1 U10461 ( .A1(n17133), .A2(\pipeline/RegFile_DEC_WB/RegBank[13][9] ), 
        .B1(n17392), .B2(\pipeline/RegFile_DEC_WB/RegBank[4][9] ), .ZN(n16123)
         );
  AOI22_X1 U10460 ( .A1(n17334), .A2(\pipeline/RegFile_DEC_WB/RegBank[10][9] ), 
        .B1(n17144), .B2(\pipeline/RegFile_DEC_WB/RegBank[3][9] ), .ZN(n16124)
         );
  AOI22_X1 U10459 ( .A1(n17338), .A2(\pipeline/RegFile_DEC_WB/RegBank[6][9] ), 
        .B1(n17142), .B2(\pipeline/RegFile_DEC_WB/RegBank[7][9] ), .ZN(n16125)
         );
  AOI22_X1 U10458 ( .A1(n17336), .A2(\pipeline/RegFile_DEC_WB/RegBank[5][9] ), 
        .B1(n17391), .B2(\pipeline/RegFile_DEC_WB/RegBank[1][9] ), .ZN(n16126)
         );
  NAND4_X1 U10457 ( .A1(n16123), .A2(n16124), .A3(n16125), .A4(n16126), .ZN(
        n16122) );
  NOR4_X1 U10456 ( .A1(n16119), .A2(n16120), .A3(n16121), .A4(n16122), .ZN(
        n14927) );
  AOI22_X1 U10455 ( .A1(n17137), .A2(\pipeline/RegFile_DEC_WB/RegBank[31][8] ), 
        .B1(n17138), .B2(\pipeline/RegFile_DEC_WB/RegBank[30][8] ), .ZN(n16116) );
  AOI22_X1 U10454 ( .A1(n17130), .A2(\pipeline/RegFile_DEC_WB/RegBank[29][8] ), 
        .B1(n17129), .B2(\pipeline/RegFile_DEC_WB/RegBank[28][8] ), .ZN(n16117) );
  AOI222_X1 U10453 ( .A1(n17135), .A2(\pipeline/RegFile_DEC_WB/RegBank[8][8] ), 
        .B1(n17132), .B2(\pipeline/RegFile_DEC_WB/RegBank[25][8] ), .C1(n17127), .C2(\pipeline/RegFile_DEC_WB/RegBank[24][8] ), .ZN(n16118) );
  AOI22_X1 U10452 ( .A1(n17143), .A2(\pipeline/RegFile_DEC_WB/RegBank[27][8] ), 
        .B1(n17145), .B2(\pipeline/RegFile_DEC_WB/RegBank[26][8] ), .ZN(n16112) );
  AOI22_X1 U10451 ( .A1(n17146), .A2(\pipeline/RegFile_DEC_WB/RegBank[23][8] ), 
        .B1(n17147), .B2(\pipeline/RegFile_DEC_WB/RegBank[22][8] ), .ZN(n16113) );
  AOI22_X1 U10450 ( .A1(n17148), .A2(\pipeline/RegFile_DEC_WB/RegBank[21][8] ), 
        .B1(n17131), .B2(\pipeline/RegFile_DEC_WB/RegBank[20][8] ), .ZN(n16114) );
  AOI22_X1 U10449 ( .A1(n17128), .A2(\pipeline/RegFile_DEC_WB/RegBank[19][8] ), 
        .B1(n17134), .B2(\pipeline/RegFile_DEC_WB/RegBank[18][8] ), .ZN(n16115) );
  NAND4_X1 U10448 ( .A1(n16112), .A2(n16113), .A3(n16114), .A4(n16115), .ZN(
        n16101) );
  AOI22_X1 U10447 ( .A1(n17141), .A2(\pipeline/RegFile_DEC_WB/RegBank[17][8] ), 
        .B1(n17341), .B2(\pipeline/RegFile_DEC_WB/RegBank[16][8] ), .ZN(n16108) );
  AOI22_X1 U10446 ( .A1(n17388), .A2(\pipeline/RegFile_DEC_WB/RegBank[9][8] ), 
        .B1(n17139), .B2(\pipeline/RegFile_DEC_WB/RegBank[2][8] ), .ZN(n16109)
         );
  AOI22_X1 U10445 ( .A1(n17136), .A2(\pipeline/RegFile_DEC_WB/RegBank[12][8] ), 
        .B1(n17389), .B2(\pipeline/RegFile_DEC_WB/RegBank[11][8] ), .ZN(n16110) );
  AOI22_X1 U10444 ( .A1(n17140), .A2(\pipeline/RegFile_DEC_WB/RegBank[14][8] ), 
        .B1(n17390), .B2(\pipeline/RegFile_DEC_WB/RegBank[15][8] ), .ZN(n16111) );
  NAND4_X1 U10443 ( .A1(n16108), .A2(n16109), .A3(n16110), .A4(n16111), .ZN(
        n16102) );
  AOI22_X1 U10442 ( .A1(n17133), .A2(\pipeline/RegFile_DEC_WB/RegBank[13][8] ), 
        .B1(n17392), .B2(\pipeline/RegFile_DEC_WB/RegBank[4][8] ), .ZN(n16104)
         );
  AOI22_X1 U10441 ( .A1(n17334), .A2(\pipeline/RegFile_DEC_WB/RegBank[10][8] ), 
        .B1(n17144), .B2(\pipeline/RegFile_DEC_WB/RegBank[3][8] ), .ZN(n16105)
         );
  AOI22_X1 U10440 ( .A1(n17338), .A2(\pipeline/RegFile_DEC_WB/RegBank[6][8] ), 
        .B1(n17142), .B2(\pipeline/RegFile_DEC_WB/RegBank[7][8] ), .ZN(n16106)
         );
  AOI22_X1 U10439 ( .A1(n17336), .A2(\pipeline/RegFile_DEC_WB/RegBank[5][8] ), 
        .B1(n17391), .B2(\pipeline/RegFile_DEC_WB/RegBank[1][8] ), .ZN(n16107)
         );
  NAND4_X1 U10438 ( .A1(n16104), .A2(n16105), .A3(n16106), .A4(n16107), .ZN(
        n16103) );
  NOR4_X1 U10437 ( .A1(n16100), .A2(n16101), .A3(n16102), .A4(n16103), .ZN(
        n14929) );
  AOI22_X1 U10436 ( .A1(n17137), .A2(\pipeline/RegFile_DEC_WB/RegBank[31][7] ), 
        .B1(n17138), .B2(\pipeline/RegFile_DEC_WB/RegBank[30][7] ), .ZN(n16097) );
  AOI22_X1 U10435 ( .A1(n17130), .A2(\pipeline/RegFile_DEC_WB/RegBank[29][7] ), 
        .B1(n17129), .B2(\pipeline/RegFile_DEC_WB/RegBank[28][7] ), .ZN(n16098) );
  AOI222_X1 U10434 ( .A1(n17135), .A2(\pipeline/RegFile_DEC_WB/RegBank[8][7] ), 
        .B1(n17132), .B2(\pipeline/RegFile_DEC_WB/RegBank[25][7] ), .C1(n17127), .C2(\pipeline/RegFile_DEC_WB/RegBank[24][7] ), .ZN(n16099) );
  AOI22_X1 U10433 ( .A1(n17143), .A2(\pipeline/RegFile_DEC_WB/RegBank[27][7] ), 
        .B1(n17145), .B2(\pipeline/RegFile_DEC_WB/RegBank[26][7] ), .ZN(n16093) );
  AOI22_X1 U10432 ( .A1(n17146), .A2(\pipeline/RegFile_DEC_WB/RegBank[23][7] ), 
        .B1(n17147), .B2(\pipeline/RegFile_DEC_WB/RegBank[22][7] ), .ZN(n16094) );
  AOI22_X1 U10431 ( .A1(n17148), .A2(\pipeline/RegFile_DEC_WB/RegBank[21][7] ), 
        .B1(n17131), .B2(\pipeline/RegFile_DEC_WB/RegBank[20][7] ), .ZN(n16095) );
  AOI22_X1 U10430 ( .A1(n17128), .A2(\pipeline/RegFile_DEC_WB/RegBank[19][7] ), 
        .B1(n17134), .B2(\pipeline/RegFile_DEC_WB/RegBank[18][7] ), .ZN(n16096) );
  NAND4_X1 U10429 ( .A1(n16093), .A2(n16094), .A3(n16095), .A4(n16096), .ZN(
        n16082) );
  AOI22_X1 U10428 ( .A1(n17141), .A2(\pipeline/RegFile_DEC_WB/RegBank[17][7] ), 
        .B1(n17341), .B2(\pipeline/RegFile_DEC_WB/RegBank[16][7] ), .ZN(n16089) );
  AOI22_X1 U10427 ( .A1(n17388), .A2(\pipeline/RegFile_DEC_WB/RegBank[9][7] ), 
        .B1(n17139), .B2(\pipeline/RegFile_DEC_WB/RegBank[2][7] ), .ZN(n16090)
         );
  AOI22_X1 U10426 ( .A1(n17136), .A2(\pipeline/RegFile_DEC_WB/RegBank[12][7] ), 
        .B1(n17389), .B2(\pipeline/RegFile_DEC_WB/RegBank[11][7] ), .ZN(n16091) );
  AOI22_X1 U10425 ( .A1(n17140), .A2(\pipeline/RegFile_DEC_WB/RegBank[14][7] ), 
        .B1(n17390), .B2(\pipeline/RegFile_DEC_WB/RegBank[15][7] ), .ZN(n16092) );
  NAND4_X1 U10424 ( .A1(n16089), .A2(n16090), .A3(n16091), .A4(n16092), .ZN(
        n16083) );
  AOI22_X1 U10423 ( .A1(n17133), .A2(\pipeline/RegFile_DEC_WB/RegBank[13][7] ), 
        .B1(n17392), .B2(\pipeline/RegFile_DEC_WB/RegBank[4][7] ), .ZN(n16085)
         );
  AOI22_X1 U10422 ( .A1(n17334), .A2(\pipeline/RegFile_DEC_WB/RegBank[10][7] ), 
        .B1(n17144), .B2(\pipeline/RegFile_DEC_WB/RegBank[3][7] ), .ZN(n16086)
         );
  AOI22_X1 U10421 ( .A1(n17338), .A2(\pipeline/RegFile_DEC_WB/RegBank[6][7] ), 
        .B1(n17142), .B2(\pipeline/RegFile_DEC_WB/RegBank[7][7] ), .ZN(n16087)
         );
  AOI22_X1 U10420 ( .A1(n17336), .A2(\pipeline/RegFile_DEC_WB/RegBank[5][7] ), 
        .B1(n17391), .B2(\pipeline/RegFile_DEC_WB/RegBank[1][7] ), .ZN(n16088)
         );
  NAND4_X1 U10419 ( .A1(n16085), .A2(n16086), .A3(n16087), .A4(n16088), .ZN(
        n16084) );
  NOR4_X1 U10418 ( .A1(n16081), .A2(n16082), .A3(n16083), .A4(n16084), .ZN(
        n14931) );
  NAND4_X1 U10417 ( .A1(n14925), .A2(n14927), .A3(n14929), .A4(n14931), .ZN(
        n16003) );
  AOI22_X1 U10416 ( .A1(n15940), .A2(\pipeline/RegFile_DEC_WB/RegBank[31][14] ), .B1(n15941), .B2(\pipeline/RegFile_DEC_WB/RegBank[30][14] ), .ZN(n16078) );
  AOI22_X1 U10415 ( .A1(n15938), .A2(\pipeline/RegFile_DEC_WB/RegBank[29][14] ), .B1(n15939), .B2(\pipeline/RegFile_DEC_WB/RegBank[28][14] ), .ZN(n16079) );
  AOI222_X1 U10414 ( .A1(n15935), .A2(\pipeline/RegFile_DEC_WB/RegBank[8][14] ), .B1(n15936), .B2(\pipeline/RegFile_DEC_WB/RegBank[25][14] ), .C1(n15937), 
        .C2(\pipeline/RegFile_DEC_WB/RegBank[24][14] ), .ZN(n16080) );
  AOI22_X1 U10413 ( .A1(n15930), .A2(\pipeline/RegFile_DEC_WB/RegBank[27][14] ), .B1(n15931), .B2(\pipeline/RegFile_DEC_WB/RegBank[26][14] ), .ZN(n16074) );
  AOI22_X1 U10412 ( .A1(n15928), .A2(\pipeline/RegFile_DEC_WB/RegBank[23][14] ), .B1(n15929), .B2(\pipeline/RegFile_DEC_WB/RegBank[22][14] ), .ZN(n16075) );
  AOI22_X1 U10411 ( .A1(n15926), .A2(\pipeline/RegFile_DEC_WB/RegBank[21][14] ), .B1(n15927), .B2(\pipeline/RegFile_DEC_WB/RegBank[20][14] ), .ZN(n16076) );
  AOI22_X1 U10410 ( .A1(n15924), .A2(\pipeline/RegFile_DEC_WB/RegBank[19][14] ), .B1(n15925), .B2(\pipeline/RegFile_DEC_WB/RegBank[18][14] ), .ZN(n16077) );
  NAND4_X1 U10409 ( .A1(n16074), .A2(n16075), .A3(n16076), .A4(n16077), .ZN(
        n16063) );
  AOI22_X1 U10408 ( .A1(n15918), .A2(\pipeline/RegFile_DEC_WB/RegBank[17][14] ), .B1(n17341), .B2(\pipeline/RegFile_DEC_WB/RegBank[16][14] ), .ZN(n16070) );
  AOI22_X1 U10407 ( .A1(n17388), .A2(\pipeline/RegFile_DEC_WB/RegBank[9][14] ), 
        .B1(n15917), .B2(\pipeline/RegFile_DEC_WB/RegBank[2][14] ), .ZN(n16071) );
  AOI22_X1 U10406 ( .A1(n15914), .A2(\pipeline/RegFile_DEC_WB/RegBank[12][14] ), .B1(n17389), .B2(\pipeline/RegFile_DEC_WB/RegBank[11][14] ), .ZN(n16072) );
  AOI22_X1 U10405 ( .A1(n15912), .A2(\pipeline/RegFile_DEC_WB/RegBank[14][14] ), .B1(n17390), .B2(\pipeline/RegFile_DEC_WB/RegBank[15][14] ), .ZN(n16073) );
  NAND4_X1 U10404 ( .A1(n16070), .A2(n16071), .A3(n16072), .A4(n16073), .ZN(
        n16064) );
  AOI22_X1 U10403 ( .A1(n15906), .A2(\pipeline/RegFile_DEC_WB/RegBank[13][14] ), .B1(n17392), .B2(\pipeline/RegFile_DEC_WB/RegBank[4][14] ), .ZN(n16066) );
  AOI22_X1 U10402 ( .A1(n17334), .A2(\pipeline/RegFile_DEC_WB/RegBank[10][14] ), .B1(n15905), .B2(\pipeline/RegFile_DEC_WB/RegBank[3][14] ), .ZN(n16067) );
  AOI22_X1 U10401 ( .A1(n17338), .A2(\pipeline/RegFile_DEC_WB/RegBank[6][14] ), 
        .B1(n15903), .B2(\pipeline/RegFile_DEC_WB/RegBank[7][14] ), .ZN(n16068) );
  AOI22_X1 U10400 ( .A1(n17336), .A2(\pipeline/RegFile_DEC_WB/RegBank[5][14] ), 
        .B1(n17391), .B2(\pipeline/RegFile_DEC_WB/RegBank[1][14] ), .ZN(n16069) );
  NAND4_X1 U10399 ( .A1(n16066), .A2(n16067), .A3(n16068), .A4(n16069), .ZN(
        n16065) );
  NOR4_X1 U10398 ( .A1(n16062), .A2(n16063), .A3(n16064), .A4(n16065), .ZN(
        n14917) );
  AOI22_X1 U10397 ( .A1(n17137), .A2(\pipeline/RegFile_DEC_WB/RegBank[31][13] ), .B1(n17138), .B2(\pipeline/RegFile_DEC_WB/RegBank[30][13] ), .ZN(n16059) );
  AOI22_X1 U10396 ( .A1(n17130), .A2(\pipeline/RegFile_DEC_WB/RegBank[29][13] ), .B1(n17129), .B2(\pipeline/RegFile_DEC_WB/RegBank[28][13] ), .ZN(n16060) );
  AOI222_X1 U10395 ( .A1(n17135), .A2(\pipeline/RegFile_DEC_WB/RegBank[8][13] ), .B1(n17132), .B2(\pipeline/RegFile_DEC_WB/RegBank[25][13] ), .C1(n17127), 
        .C2(\pipeline/RegFile_DEC_WB/RegBank[24][13] ), .ZN(n16061) );
  AOI22_X1 U10394 ( .A1(n17143), .A2(\pipeline/RegFile_DEC_WB/RegBank[27][13] ), .B1(n17145), .B2(\pipeline/RegFile_DEC_WB/RegBank[26][13] ), .ZN(n16055) );
  AOI22_X1 U10393 ( .A1(n17146), .A2(\pipeline/RegFile_DEC_WB/RegBank[23][13] ), .B1(n17147), .B2(\pipeline/RegFile_DEC_WB/RegBank[22][13] ), .ZN(n16056) );
  AOI22_X1 U10392 ( .A1(n17148), .A2(\pipeline/RegFile_DEC_WB/RegBank[21][13] ), .B1(n17131), .B2(\pipeline/RegFile_DEC_WB/RegBank[20][13] ), .ZN(n16057) );
  AOI22_X1 U10391 ( .A1(n17128), .A2(\pipeline/RegFile_DEC_WB/RegBank[19][13] ), .B1(n17134), .B2(\pipeline/RegFile_DEC_WB/RegBank[18][13] ), .ZN(n16058) );
  NAND4_X1 U10390 ( .A1(n16055), .A2(n16056), .A3(n16057), .A4(n16058), .ZN(
        n16044) );
  AOI22_X1 U10389 ( .A1(n17141), .A2(\pipeline/RegFile_DEC_WB/RegBank[17][13] ), .B1(n17341), .B2(\pipeline/RegFile_DEC_WB/RegBank[16][13] ), .ZN(n16051) );
  AOI22_X1 U10388 ( .A1(n17388), .A2(\pipeline/RegFile_DEC_WB/RegBank[9][13] ), 
        .B1(n17139), .B2(\pipeline/RegFile_DEC_WB/RegBank[2][13] ), .ZN(n16052) );
  AOI22_X1 U10387 ( .A1(n17136), .A2(\pipeline/RegFile_DEC_WB/RegBank[12][13] ), .B1(n17389), .B2(\pipeline/RegFile_DEC_WB/RegBank[11][13] ), .ZN(n16053) );
  AOI22_X1 U10386 ( .A1(n17140), .A2(\pipeline/RegFile_DEC_WB/RegBank[14][13] ), .B1(n17390), .B2(\pipeline/RegFile_DEC_WB/RegBank[15][13] ), .ZN(n16054) );
  NAND4_X1 U10385 ( .A1(n16051), .A2(n16052), .A3(n16053), .A4(n16054), .ZN(
        n16045) );
  AOI22_X1 U10384 ( .A1(n17133), .A2(\pipeline/RegFile_DEC_WB/RegBank[13][13] ), .B1(n17392), .B2(\pipeline/RegFile_DEC_WB/RegBank[4][13] ), .ZN(n16047) );
  AOI22_X1 U10383 ( .A1(n17334), .A2(\pipeline/RegFile_DEC_WB/RegBank[10][13] ), .B1(n17144), .B2(\pipeline/RegFile_DEC_WB/RegBank[3][13] ), .ZN(n16048) );
  AOI22_X1 U10382 ( .A1(n17338), .A2(\pipeline/RegFile_DEC_WB/RegBank[6][13] ), 
        .B1(n17142), .B2(\pipeline/RegFile_DEC_WB/RegBank[7][13] ), .ZN(n16049) );
  AOI22_X1 U10381 ( .A1(n17336), .A2(\pipeline/RegFile_DEC_WB/RegBank[5][13] ), 
        .B1(n17391), .B2(\pipeline/RegFile_DEC_WB/RegBank[1][13] ), .ZN(n16050) );
  NAND4_X1 U10380 ( .A1(n16047), .A2(n16048), .A3(n16049), .A4(n16050), .ZN(
        n16046) );
  NOR4_X1 U10379 ( .A1(n16043), .A2(n16044), .A3(n16045), .A4(n16046), .ZN(
        n14919) );
  AOI22_X1 U10378 ( .A1(n17137), .A2(\pipeline/RegFile_DEC_WB/RegBank[31][12] ), .B1(n17138), .B2(\pipeline/RegFile_DEC_WB/RegBank[30][12] ), .ZN(n16040) );
  AOI22_X1 U10377 ( .A1(n17130), .A2(\pipeline/RegFile_DEC_WB/RegBank[29][12] ), .B1(n17129), .B2(\pipeline/RegFile_DEC_WB/RegBank[28][12] ), .ZN(n16041) );
  AOI222_X1 U10376 ( .A1(n17135), .A2(\pipeline/RegFile_DEC_WB/RegBank[8][12] ), .B1(n17132), .B2(\pipeline/RegFile_DEC_WB/RegBank[25][12] ), .C1(n17127), 
        .C2(\pipeline/RegFile_DEC_WB/RegBank[24][12] ), .ZN(n16042) );
  AOI22_X1 U10375 ( .A1(n17143), .A2(\pipeline/RegFile_DEC_WB/RegBank[27][12] ), .B1(n17145), .B2(\pipeline/RegFile_DEC_WB/RegBank[26][12] ), .ZN(n16036) );
  AOI22_X1 U10374 ( .A1(n17146), .A2(\pipeline/RegFile_DEC_WB/RegBank[23][12] ), .B1(n17147), .B2(\pipeline/RegFile_DEC_WB/RegBank[22][12] ), .ZN(n16037) );
  AOI22_X1 U10373 ( .A1(n17148), .A2(\pipeline/RegFile_DEC_WB/RegBank[21][12] ), .B1(n17131), .B2(\pipeline/RegFile_DEC_WB/RegBank[20][12] ), .ZN(n16038) );
  AOI22_X1 U10372 ( .A1(n17128), .A2(\pipeline/RegFile_DEC_WB/RegBank[19][12] ), .B1(n17134), .B2(\pipeline/RegFile_DEC_WB/RegBank[18][12] ), .ZN(n16039) );
  NAND4_X1 U10371 ( .A1(n16036), .A2(n16037), .A3(n16038), .A4(n16039), .ZN(
        n16025) );
  AOI22_X1 U10370 ( .A1(n17141), .A2(\pipeline/RegFile_DEC_WB/RegBank[17][12] ), .B1(n17341), .B2(\pipeline/RegFile_DEC_WB/RegBank[16][12] ), .ZN(n16032) );
  AOI22_X1 U10369 ( .A1(n17388), .A2(\pipeline/RegFile_DEC_WB/RegBank[9][12] ), 
        .B1(n17139), .B2(\pipeline/RegFile_DEC_WB/RegBank[2][12] ), .ZN(n16033) );
  AOI22_X1 U10368 ( .A1(n17136), .A2(\pipeline/RegFile_DEC_WB/RegBank[12][12] ), .B1(n17389), .B2(\pipeline/RegFile_DEC_WB/RegBank[11][12] ), .ZN(n16034) );
  AOI22_X1 U10367 ( .A1(n17140), .A2(\pipeline/RegFile_DEC_WB/RegBank[14][12] ), .B1(n17390), .B2(\pipeline/RegFile_DEC_WB/RegBank[15][12] ), .ZN(n16035) );
  NAND4_X1 U10366 ( .A1(n16032), .A2(n16033), .A3(n16034), .A4(n16035), .ZN(
        n16026) );
  AOI22_X1 U10365 ( .A1(n17133), .A2(\pipeline/RegFile_DEC_WB/RegBank[13][12] ), .B1(n17392), .B2(\pipeline/RegFile_DEC_WB/RegBank[4][12] ), .ZN(n16028) );
  AOI22_X1 U10364 ( .A1(n17334), .A2(\pipeline/RegFile_DEC_WB/RegBank[10][12] ), .B1(n17144), .B2(\pipeline/RegFile_DEC_WB/RegBank[3][12] ), .ZN(n16029) );
  AOI22_X1 U10363 ( .A1(n17338), .A2(\pipeline/RegFile_DEC_WB/RegBank[6][12] ), 
        .B1(n17142), .B2(\pipeline/RegFile_DEC_WB/RegBank[7][12] ), .ZN(n16030) );
  AOI22_X1 U10362 ( .A1(n17336), .A2(\pipeline/RegFile_DEC_WB/RegBank[5][12] ), 
        .B1(n17391), .B2(\pipeline/RegFile_DEC_WB/RegBank[1][12] ), .ZN(n16031) );
  NAND4_X1 U10361 ( .A1(n16028), .A2(n16029), .A3(n16030), .A4(n16031), .ZN(
        n16027) );
  NOR4_X1 U10360 ( .A1(n16024), .A2(n16025), .A3(n16026), .A4(n16027), .ZN(
        n14921) );
  AOI22_X1 U10359 ( .A1(n17137), .A2(\pipeline/RegFile_DEC_WB/RegBank[31][11] ), .B1(n17138), .B2(\pipeline/RegFile_DEC_WB/RegBank[30][11] ), .ZN(n16021) );
  AOI22_X1 U10358 ( .A1(n17130), .A2(\pipeline/RegFile_DEC_WB/RegBank[29][11] ), .B1(n17129), .B2(\pipeline/RegFile_DEC_WB/RegBank[28][11] ), .ZN(n16022) );
  AOI222_X1 U10357 ( .A1(n17135), .A2(\pipeline/RegFile_DEC_WB/RegBank[8][11] ), .B1(n17132), .B2(\pipeline/RegFile_DEC_WB/RegBank[25][11] ), .C1(n17127), 
        .C2(\pipeline/RegFile_DEC_WB/RegBank[24][11] ), .ZN(n16023) );
  AOI22_X1 U10356 ( .A1(n17143), .A2(\pipeline/RegFile_DEC_WB/RegBank[27][11] ), .B1(n17145), .B2(\pipeline/RegFile_DEC_WB/RegBank[26][11] ), .ZN(n16017) );
  AOI22_X1 U10355 ( .A1(n17146), .A2(\pipeline/RegFile_DEC_WB/RegBank[23][11] ), .B1(n17147), .B2(\pipeline/RegFile_DEC_WB/RegBank[22][11] ), .ZN(n16018) );
  AOI22_X1 U10354 ( .A1(n17148), .A2(\pipeline/RegFile_DEC_WB/RegBank[21][11] ), .B1(n17131), .B2(\pipeline/RegFile_DEC_WB/RegBank[20][11] ), .ZN(n16019) );
  AOI22_X1 U10353 ( .A1(n17128), .A2(\pipeline/RegFile_DEC_WB/RegBank[19][11] ), .B1(n17134), .B2(\pipeline/RegFile_DEC_WB/RegBank[18][11] ), .ZN(n16020) );
  NAND4_X1 U10352 ( .A1(n16017), .A2(n16018), .A3(n16019), .A4(n16020), .ZN(
        n16006) );
  AOI22_X1 U10351 ( .A1(n17141), .A2(\pipeline/RegFile_DEC_WB/RegBank[17][11] ), .B1(n17342), .B2(\pipeline/RegFile_DEC_WB/RegBank[16][11] ), .ZN(n16013) );
  AOI22_X1 U10350 ( .A1(n17388), .A2(\pipeline/RegFile_DEC_WB/RegBank[9][11] ), 
        .B1(n17139), .B2(\pipeline/RegFile_DEC_WB/RegBank[2][11] ), .ZN(n16014) );
  AOI22_X1 U10349 ( .A1(n17136), .A2(\pipeline/RegFile_DEC_WB/RegBank[12][11] ), .B1(n17389), .B2(\pipeline/RegFile_DEC_WB/RegBank[11][11] ), .ZN(n16015) );
  AOI22_X1 U10348 ( .A1(n17140), .A2(\pipeline/RegFile_DEC_WB/RegBank[14][11] ), .B1(n17390), .B2(\pipeline/RegFile_DEC_WB/RegBank[15][11] ), .ZN(n16016) );
  NAND4_X1 U10347 ( .A1(n16013), .A2(n16014), .A3(n16015), .A4(n16016), .ZN(
        n16007) );
  AOI22_X1 U10346 ( .A1(n17133), .A2(\pipeline/RegFile_DEC_WB/RegBank[13][11] ), .B1(n17392), .B2(\pipeline/RegFile_DEC_WB/RegBank[4][11] ), .ZN(n16009) );
  AOI22_X1 U10345 ( .A1(n17335), .A2(\pipeline/RegFile_DEC_WB/RegBank[10][11] ), .B1(n17144), .B2(\pipeline/RegFile_DEC_WB/RegBank[3][11] ), .ZN(n16010) );
  AOI22_X1 U10344 ( .A1(n17339), .A2(\pipeline/RegFile_DEC_WB/RegBank[6][11] ), 
        .B1(n17142), .B2(\pipeline/RegFile_DEC_WB/RegBank[7][11] ), .ZN(n16011) );
  AOI22_X1 U10343 ( .A1(n17337), .A2(\pipeline/RegFile_DEC_WB/RegBank[5][11] ), 
        .B1(n17391), .B2(\pipeline/RegFile_DEC_WB/RegBank[1][11] ), .ZN(n16012) );
  NAND4_X1 U10342 ( .A1(n16009), .A2(n16010), .A3(n16011), .A4(n16012), .ZN(
        n16008) );
  NOR4_X1 U10341 ( .A1(n16005), .A2(n16006), .A3(n16007), .A4(n16008), .ZN(
        n14923) );
  NAND4_X1 U10340 ( .A1(n14917), .A2(n14919), .A3(n14921), .A4(n14923), .ZN(
        n16004) );
  NOR4_X1 U10339 ( .A1(n16001), .A2(n16002), .A3(n16003), .A4(n16004), .ZN(
        n16000) );
  NAND4_X1 U10338 ( .A1(n14933), .A2(n14935), .A3(n15999), .A4(n16000), .ZN(
        n15890) );
  AOI22_X1 U10337 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[31][30] ), .A2(n17137), .B1(\pipeline/RegFile_DEC_WB/RegBank[30][30] ), .B2(n17138), .ZN(n15996) );
  AOI22_X1 U10336 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[29][30] ), .A2(n17130), .B1(\pipeline/RegFile_DEC_WB/RegBank[28][30] ), .B2(n17129), .ZN(n15997) );
  AOI222_X1 U10335 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[8][30] ), .A2(n17135), .B1(\pipeline/RegFile_DEC_WB/RegBank[25][30] ), .B2(n17132), .C1(
        \pipeline/RegFile_DEC_WB/RegBank[24][30] ), .C2(n17127), .ZN(n15998)
         );
  AOI22_X1 U10334 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[27][30] ), .A2(n17143), .B1(\pipeline/RegFile_DEC_WB/RegBank[26][30] ), .B2(n17145), .ZN(n15992) );
  AOI22_X1 U10333 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[23][30] ), .A2(n17146), .B1(\pipeline/RegFile_DEC_WB/RegBank[22][30] ), .B2(n17147), .ZN(n15993) );
  AOI22_X1 U10332 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[21][30] ), .A2(n17148), .B1(\pipeline/RegFile_DEC_WB/RegBank[20][30] ), .B2(n17131), .ZN(n15994) );
  AOI22_X1 U10331 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[19][30] ), .A2(n17128), .B1(\pipeline/RegFile_DEC_WB/RegBank[18][30] ), .B2(n17134), .ZN(n15995) );
  NAND4_X1 U10330 ( .A1(n15992), .A2(n15993), .A3(n15994), .A4(n15995), .ZN(
        n15981) );
  AOI22_X1 U10329 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[17][30] ), .A2(n17141), .B1(\pipeline/RegFile_DEC_WB/RegBank[16][30] ), .B2(n17341), .ZN(n15988) );
  AOI22_X1 U10328 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[9][30] ), .A2(n17388), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[2][30] ), .B2(n17139), .ZN(n15989) );
  AOI22_X1 U10327 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[12][30] ), .A2(n17136), .B1(\pipeline/RegFile_DEC_WB/RegBank[11][30] ), .B2(n17389), .ZN(n15990) );
  AOI22_X1 U10326 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[14][30] ), .A2(n17140), .B1(\pipeline/RegFile_DEC_WB/RegBank[15][30] ), .B2(n17390), .ZN(n15991) );
  NAND4_X1 U10325 ( .A1(n15988), .A2(n15989), .A3(n15990), .A4(n15991), .ZN(
        n15982) );
  AOI22_X1 U10324 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[13][30] ), .A2(n17133), .B1(\pipeline/RegFile_DEC_WB/RegBank[4][30] ), .B2(n17392), .ZN(n15984) );
  AOI22_X1 U10323 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[10][30] ), .A2(n17334), .B1(\pipeline/RegFile_DEC_WB/RegBank[3][30] ), .B2(n17144), .ZN(n15985) );
  AOI22_X1 U10322 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[6][30] ), .A2(n17338), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[7][30] ), .B2(n17142), .ZN(n15986) );
  AOI22_X1 U10321 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[5][30] ), .A2(n17336), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[1][30] ), .B2(n17391), .ZN(n15987) );
  NAND4_X1 U10320 ( .A1(n15984), .A2(n15985), .A3(n15986), .A4(n15987), .ZN(
        n15983) );
  NOR4_X1 U10319 ( .A1(n15980), .A2(n15981), .A3(n15982), .A4(n15983), .ZN(
        n14885) );
  AOI22_X1 U10318 ( .A1(n15940), .A2(\pipeline/RegFile_DEC_WB/RegBank[31][29] ), .B1(n15941), .B2(\pipeline/RegFile_DEC_WB/RegBank[30][29] ), .ZN(n15977) );
  AOI22_X1 U10317 ( .A1(n15938), .A2(\pipeline/RegFile_DEC_WB/RegBank[29][29] ), .B1(n15939), .B2(\pipeline/RegFile_DEC_WB/RegBank[28][29] ), .ZN(n15978) );
  AOI222_X1 U10316 ( .A1(n15935), .A2(\pipeline/RegFile_DEC_WB/RegBank[8][29] ), .B1(n15936), .B2(\pipeline/RegFile_DEC_WB/RegBank[25][29] ), .C1(n15937), 
        .C2(\pipeline/RegFile_DEC_WB/RegBank[24][29] ), .ZN(n15979) );
  AOI22_X1 U10315 ( .A1(n15930), .A2(\pipeline/RegFile_DEC_WB/RegBank[27][29] ), .B1(n15931), .B2(\pipeline/RegFile_DEC_WB/RegBank[26][29] ), .ZN(n15973) );
  AOI22_X1 U10314 ( .A1(n15928), .A2(\pipeline/RegFile_DEC_WB/RegBank[23][29] ), .B1(n15929), .B2(\pipeline/RegFile_DEC_WB/RegBank[22][29] ), .ZN(n15974) );
  AOI22_X1 U10313 ( .A1(n15926), .A2(\pipeline/RegFile_DEC_WB/RegBank[21][29] ), .B1(n15927), .B2(\pipeline/RegFile_DEC_WB/RegBank[20][29] ), .ZN(n15975) );
  AOI22_X1 U10312 ( .A1(n15924), .A2(\pipeline/RegFile_DEC_WB/RegBank[19][29] ), .B1(n15925), .B2(\pipeline/RegFile_DEC_WB/RegBank[18][29] ), .ZN(n15976) );
  NAND4_X1 U10311 ( .A1(n15973), .A2(n15974), .A3(n15975), .A4(n15976), .ZN(
        n15962) );
  AOI22_X1 U10310 ( .A1(n15918), .A2(\pipeline/RegFile_DEC_WB/RegBank[17][29] ), .B1(n17342), .B2(\pipeline/RegFile_DEC_WB/RegBank[16][29] ), .ZN(n15969) );
  AOI22_X1 U10309 ( .A1(n17388), .A2(\pipeline/RegFile_DEC_WB/RegBank[9][29] ), 
        .B1(n15917), .B2(\pipeline/RegFile_DEC_WB/RegBank[2][29] ), .ZN(n15970) );
  AOI22_X1 U10308 ( .A1(n15914), .A2(\pipeline/RegFile_DEC_WB/RegBank[12][29] ), .B1(n17389), .B2(\pipeline/RegFile_DEC_WB/RegBank[11][29] ), .ZN(n15971) );
  AOI22_X1 U10307 ( .A1(n15912), .A2(\pipeline/RegFile_DEC_WB/RegBank[14][29] ), .B1(n17390), .B2(\pipeline/RegFile_DEC_WB/RegBank[15][29] ), .ZN(n15972) );
  NAND4_X1 U10306 ( .A1(n15969), .A2(n15970), .A3(n15971), .A4(n15972), .ZN(
        n15963) );
  AOI22_X1 U10305 ( .A1(n15906), .A2(\pipeline/RegFile_DEC_WB/RegBank[13][29] ), .B1(n17392), .B2(\pipeline/RegFile_DEC_WB/RegBank[4][29] ), .ZN(n15965) );
  AOI22_X1 U10304 ( .A1(n17335), .A2(\pipeline/RegFile_DEC_WB/RegBank[10][29] ), .B1(n15905), .B2(\pipeline/RegFile_DEC_WB/RegBank[3][29] ), .ZN(n15966) );
  AOI22_X1 U10303 ( .A1(n17339), .A2(\pipeline/RegFile_DEC_WB/RegBank[6][29] ), 
        .B1(n15903), .B2(\pipeline/RegFile_DEC_WB/RegBank[7][29] ), .ZN(n15967) );
  AOI22_X1 U10302 ( .A1(n17337), .A2(\pipeline/RegFile_DEC_WB/RegBank[5][29] ), 
        .B1(n17391), .B2(\pipeline/RegFile_DEC_WB/RegBank[1][29] ), .ZN(n15968) );
  NAND4_X1 U10301 ( .A1(n15965), .A2(n15966), .A3(n15967), .A4(n15968), .ZN(
        n15964) );
  NOR4_X1 U10300 ( .A1(n15961), .A2(n15962), .A3(n15963), .A4(n15964), .ZN(
        n14887) );
  AOI22_X1 U10299 ( .A1(n17137), .A2(\pipeline/RegFile_DEC_WB/RegBank[31][28] ), .B1(n17138), .B2(\pipeline/RegFile_DEC_WB/RegBank[30][28] ), .ZN(n15958) );
  AOI22_X1 U10298 ( .A1(n17130), .A2(\pipeline/RegFile_DEC_WB/RegBank[29][28] ), .B1(n17129), .B2(\pipeline/RegFile_DEC_WB/RegBank[28][28] ), .ZN(n15959) );
  AOI222_X1 U10297 ( .A1(n17135), .A2(\pipeline/RegFile_DEC_WB/RegBank[8][28] ), .B1(n17132), .B2(\pipeline/RegFile_DEC_WB/RegBank[25][28] ), .C1(n17127), 
        .C2(\pipeline/RegFile_DEC_WB/RegBank[24][28] ), .ZN(n15960) );
  AOI22_X1 U10296 ( .A1(n17143), .A2(\pipeline/RegFile_DEC_WB/RegBank[27][28] ), .B1(n17145), .B2(\pipeline/RegFile_DEC_WB/RegBank[26][28] ), .ZN(n15954) );
  AOI22_X1 U10295 ( .A1(n17146), .A2(\pipeline/RegFile_DEC_WB/RegBank[23][28] ), .B1(n17147), .B2(\pipeline/RegFile_DEC_WB/RegBank[22][28] ), .ZN(n15955) );
  AOI22_X1 U10294 ( .A1(n17148), .A2(\pipeline/RegFile_DEC_WB/RegBank[21][28] ), .B1(n17131), .B2(\pipeline/RegFile_DEC_WB/RegBank[20][28] ), .ZN(n15956) );
  AOI22_X1 U10293 ( .A1(n17128), .A2(\pipeline/RegFile_DEC_WB/RegBank[19][28] ), .B1(n17134), .B2(\pipeline/RegFile_DEC_WB/RegBank[18][28] ), .ZN(n15957) );
  NAND4_X1 U10292 ( .A1(n15954), .A2(n15955), .A3(n15956), .A4(n15957), .ZN(
        n15943) );
  AOI22_X1 U10291 ( .A1(n17141), .A2(\pipeline/RegFile_DEC_WB/RegBank[17][28] ), .B1(n17342), .B2(\pipeline/RegFile_DEC_WB/RegBank[16][28] ), .ZN(n15950) );
  AOI22_X1 U10290 ( .A1(n17388), .A2(\pipeline/RegFile_DEC_WB/RegBank[9][28] ), 
        .B1(n17139), .B2(\pipeline/RegFile_DEC_WB/RegBank[2][28] ), .ZN(n15951) );
  AOI22_X1 U10289 ( .A1(n17136), .A2(\pipeline/RegFile_DEC_WB/RegBank[12][28] ), .B1(n17389), .B2(\pipeline/RegFile_DEC_WB/RegBank[11][28] ), .ZN(n15952) );
  AOI22_X1 U10288 ( .A1(n17140), .A2(\pipeline/RegFile_DEC_WB/RegBank[14][28] ), .B1(n17390), .B2(\pipeline/RegFile_DEC_WB/RegBank[15][28] ), .ZN(n15953) );
  NAND4_X1 U10287 ( .A1(n15950), .A2(n15951), .A3(n15952), .A4(n15953), .ZN(
        n15944) );
  AOI22_X1 U10286 ( .A1(n17133), .A2(\pipeline/RegFile_DEC_WB/RegBank[13][28] ), .B1(n17392), .B2(\pipeline/RegFile_DEC_WB/RegBank[4][28] ), .ZN(n15946) );
  AOI22_X1 U10285 ( .A1(n17335), .A2(\pipeline/RegFile_DEC_WB/RegBank[10][28] ), .B1(n17144), .B2(\pipeline/RegFile_DEC_WB/RegBank[3][28] ), .ZN(n15947) );
  AOI22_X1 U10284 ( .A1(n17339), .A2(\pipeline/RegFile_DEC_WB/RegBank[6][28] ), 
        .B1(n17142), .B2(\pipeline/RegFile_DEC_WB/RegBank[7][28] ), .ZN(n15948) );
  AOI22_X1 U10283 ( .A1(n17337), .A2(\pipeline/RegFile_DEC_WB/RegBank[5][28] ), 
        .B1(n17391), .B2(\pipeline/RegFile_DEC_WB/RegBank[1][28] ), .ZN(n15949) );
  NAND4_X1 U10282 ( .A1(n15946), .A2(n15947), .A3(n15948), .A4(n15949), .ZN(
        n15945) );
  NOR4_X1 U10281 ( .A1(n15942), .A2(n15943), .A3(n15944), .A4(n15945), .ZN(
        n14889) );
  AOI22_X1 U10280 ( .A1(n17137), .A2(\pipeline/RegFile_DEC_WB/RegBank[31][27] ), .B1(n17138), .B2(\pipeline/RegFile_DEC_WB/RegBank[30][27] ), .ZN(n15932) );
  AOI22_X1 U10279 ( .A1(n17130), .A2(\pipeline/RegFile_DEC_WB/RegBank[29][27] ), .B1(n17129), .B2(\pipeline/RegFile_DEC_WB/RegBank[28][27] ), .ZN(n15933) );
  AOI222_X1 U10278 ( .A1(n17135), .A2(\pipeline/RegFile_DEC_WB/RegBank[8][27] ), .B1(n17132), .B2(\pipeline/RegFile_DEC_WB/RegBank[25][27] ), .C1(n17127), 
        .C2(\pipeline/RegFile_DEC_WB/RegBank[24][27] ), .ZN(n15934) );
  AOI22_X1 U10277 ( .A1(n17143), .A2(\pipeline/RegFile_DEC_WB/RegBank[27][27] ), .B1(n17145), .B2(\pipeline/RegFile_DEC_WB/RegBank[26][27] ), .ZN(n15920) );
  AOI22_X1 U10276 ( .A1(n17146), .A2(\pipeline/RegFile_DEC_WB/RegBank[23][27] ), .B1(n17147), .B2(\pipeline/RegFile_DEC_WB/RegBank[22][27] ), .ZN(n15921) );
  AOI22_X1 U10275 ( .A1(n17148), .A2(\pipeline/RegFile_DEC_WB/RegBank[21][27] ), .B1(n17131), .B2(\pipeline/RegFile_DEC_WB/RegBank[20][27] ), .ZN(n15922) );
  AOI22_X1 U10274 ( .A1(n17128), .A2(\pipeline/RegFile_DEC_WB/RegBank[19][27] ), .B1(n17134), .B2(\pipeline/RegFile_DEC_WB/RegBank[18][27] ), .ZN(n15923) );
  NAND4_X1 U10273 ( .A1(n15920), .A2(n15921), .A3(n15922), .A4(n15923), .ZN(
        n15893) );
  AOI22_X1 U10272 ( .A1(n17141), .A2(\pipeline/RegFile_DEC_WB/RegBank[17][27] ), .B1(n17342), .B2(\pipeline/RegFile_DEC_WB/RegBank[16][27] ), .ZN(n15908) );
  AOI22_X1 U10271 ( .A1(n15916), .A2(\pipeline/RegFile_DEC_WB/RegBank[9][27] ), 
        .B1(n17139), .B2(\pipeline/RegFile_DEC_WB/RegBank[2][27] ), .ZN(n15909) );
  AOI22_X1 U10270 ( .A1(n17136), .A2(\pipeline/RegFile_DEC_WB/RegBank[12][27] ), .B1(n15915), .B2(\pipeline/RegFile_DEC_WB/RegBank[11][27] ), .ZN(n15910) );
  AOI22_X1 U10269 ( .A1(n17140), .A2(\pipeline/RegFile_DEC_WB/RegBank[14][27] ), .B1(n15913), .B2(\pipeline/RegFile_DEC_WB/RegBank[15][27] ), .ZN(n15911) );
  NAND4_X1 U10268 ( .A1(n15908), .A2(n15909), .A3(n15910), .A4(n15911), .ZN(
        n15894) );
  AOI22_X1 U10267 ( .A1(n17133), .A2(\pipeline/RegFile_DEC_WB/RegBank[13][27] ), .B1(n15907), .B2(\pipeline/RegFile_DEC_WB/RegBank[4][27] ), .ZN(n15896) );
  AOI22_X1 U10266 ( .A1(n17335), .A2(\pipeline/RegFile_DEC_WB/RegBank[10][27] ), .B1(n17144), .B2(\pipeline/RegFile_DEC_WB/RegBank[3][27] ), .ZN(n15897) );
  AOI22_X1 U10265 ( .A1(n17339), .A2(\pipeline/RegFile_DEC_WB/RegBank[6][27] ), 
        .B1(n17142), .B2(\pipeline/RegFile_DEC_WB/RegBank[7][27] ), .ZN(n15898) );
  AOI22_X1 U10264 ( .A1(n17337), .A2(\pipeline/RegFile_DEC_WB/RegBank[5][27] ), 
        .B1(n15901), .B2(\pipeline/RegFile_DEC_WB/RegBank[1][27] ), .ZN(n15899) );
  NAND4_X1 U10263 ( .A1(n15896), .A2(n15897), .A3(n15898), .A4(n15899), .ZN(
        n15895) );
  NOR4_X1 U10262 ( .A1(n15892), .A2(n15893), .A3(n15894), .A4(n15895), .ZN(
        n14891) );
  NAND4_X1 U10261 ( .A1(n14885), .A2(n14887), .A3(n14889), .A4(n14891), .ZN(
        n15891) );
  NAND4_X1 U10259 ( .A1(n17423), .A2(n17363), .A3(n17322), .A4(n17310), .ZN(
        n15866) );
  NAND4_X1 U10258 ( .A1(n17427), .A2(n17324), .A3(n17366), .A4(n17311), .ZN(
        n15867) );
  NAND4_X1 U10257 ( .A1(n17344), .A2(n17319), .A3(n17307), .A4(n17395), .ZN(
        n15868) );
  NAND4_X1 U10256 ( .A1(n17309), .A2(n17364), .A3(n17323), .A4(n17426), .ZN(
        n15869) );
  NOR4_X1 U10255 ( .A1(n15866), .A2(n15867), .A3(n15868), .A4(n15869), .ZN(
        n15844) );
  NAND4_X1 U10254 ( .A1(n17394), .A2(n17343), .A3(n17318), .A4(n17305), .ZN(
        n15846) );
  NAND4_X1 U10253 ( .A1(n17396), .A2(n17369), .A3(n17321), .A4(n17306), .ZN(
        n15847) );
  NAND4_X1 U10252 ( .A1(n17424), .A2(n17325), .A3(n17312), .A4(n17365), .ZN(
        n15848) );
  NAND4_X1 U10251 ( .A1(n17425), .A2(n17320), .A3(n17308), .A4(n17362), .ZN(
        n15849) );
  NOR4_X1 U10250 ( .A1(n15846), .A2(n15847), .A3(n15848), .A4(n15849), .ZN(
        n15845) );
  NAND2_X1 U10245 ( .A1(\pipeline/inst_IFID_DEC[26] ), .A2(n17347), .ZN(n14059) );
  NAND2_X1 U10241 ( .A1(n14126), .A2(n14167), .ZN(n15840) );
  NOR3_X1 U10238 ( .A1(n13281), .A2(n14176), .A3(n14186), .ZN(n14125) );
  XNOR2_X1 U11431 ( .A(\pipeline/regDst_to_mem[0] ), .B(
        \pipeline/Reg2_Addr_to_exe [0]), .ZN(n16789) );
  OAI221_X1 U11423 ( .B1(n17304), .B2(\pipeline/Reg2_Addr_to_exe [1]), .C1(
        n17386), .C2(\pipeline/Reg2_Addr_to_exe [4]), .A(n16784), .ZN(n16779)
         );
  NOR2_X1 U11321 ( .A1(\pipeline/EXE_controls_in_EXEcute [0]), .A2(n13877), 
        .ZN(n16731) );
  AOI22_X1 U11320 ( .A1(n16607), .A2(\pipeline/Alu_Out_Addr_to_mem[13] ), .B1(
        n17670), .B2(\pipeline/data_to_RF_from_WB[13] ), .ZN(n16732) );
  OAI21_X1 U11319 ( .B1(n17120), .B2(n16731), .A(n16732), .ZN(n16730) );
  OAI21_X1 U11318 ( .B1(\pipeline/immediate_to_exe [13]), .B2(n17327), .A(
        n16730), .ZN(n15427) );
  XNOR2_X1 U11316 ( .A(n17381), .B(n15426), .ZN(n16659) );
  XNOR2_X1 U11466 ( .A(n17645), .B(\pipeline/Reg1_Addr_to_exe [1]), .ZN(n16808) );
  NOR2_X1 U11465 ( .A1(n16808), .A2(n16809), .ZN(n16807) );
  XNOR2_X1 U11472 ( .A(n17646), .B(\pipeline/Reg1_Addr_to_exe [2]), .ZN(n16795) );
  AOI22_X1 U11314 ( .A1(n17663), .A2(\pipeline/Alu_Out_Addr_to_mem[13] ), .B1(
        n17664), .B2(n13958), .ZN(n16729) );
  NAND2_X1 U11312 ( .A1(n16659), .A2(\pipeline/stageE/input1_to_ALU [13]), 
        .ZN(n15416) );
  NAND2_X1 U11233 ( .A1(n16691), .A2(n12649), .ZN(n15053) );
  AOI22_X1 U11230 ( .A1(n17663), .A2(\pipeline/Alu_Out_Addr_to_mem[3] ), .B1(
        n17664), .B2(n13844), .ZN(n16689) );
  NOR2_X1 U11227 ( .A1(\pipeline/EXE_controls_in_EXEcute [0]), .A2(n13838), 
        .ZN(n16685) );
  AOI22_X1 U11226 ( .A1(n16607), .A2(\pipeline/Alu_Out_Addr_to_mem[4] ), .B1(
        n15123), .B2(\pipeline/data_to_RF_from_WB[4] ), .ZN(n16686) );
  NOR2_X1 U11225 ( .A1(\pipeline/immediate_to_exe [4]), .A2(n17327), .ZN(
        n16687) );
  AOI221_X1 U11224 ( .B1(n16685), .B2(n16686), .C1(n17120), .C2(n16686), .A(
        n16687), .ZN(n4376) );
  OAI22_X1 U11222 ( .A1(n17381), .A2(n17737), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .B2(
        \pipeline/stageE/EXE_ALU/add_alu/sCout[0] ), .ZN(n16683) );
  AOI22_X1 U11220 ( .A1(n17663), .A2(\pipeline/Alu_Out_Addr_to_mem[4] ), .B1(
        n17664), .B2(n13836), .ZN(n16684) );
  NAND2_X1 U11215 ( .A1(n15564), .A2(n16683), .ZN(n15568) );
  NOR2_X1 U11279 ( .A1(\pipeline/EXE_controls_in_EXEcute [0]), .A2(n13834), 
        .ZN(n16711) );
  AOI22_X1 U11278 ( .A1(n16607), .A2(\pipeline/Alu_Out_Addr_to_mem[5] ), .B1(
        n17670), .B2(\pipeline/data_to_RF_from_WB[5] ), .ZN(n16712) );
  OAI21_X1 U11277 ( .B1(n17120), .B2(n16711), .A(n16712), .ZN(n16710) );
  OAI21_X1 U11276 ( .B1(\pipeline/immediate_to_exe [5]), .B2(n17327), .A(
        n16710), .ZN(n15553) );
  NOR2_X1 U11272 ( .A1(n16677), .A2(\pipeline/stageE/input1_to_ALU [5]), .ZN(
        n15542) );
  NOR2_X1 U11213 ( .A1(\pipeline/EXE_controls_in_EXEcute [0]), .A2(n13843), 
        .ZN(n16680) );
  AOI22_X1 U11212 ( .A1(n17665), .A2(\pipeline/Alu_Out_Addr_to_mem[6] ), .B1(
        n17123), .B2(\pipeline/data_to_RF_from_WB[6] ), .ZN(n16681) );
  OAI21_X1 U11211 ( .B1(n17120), .B2(n16680), .A(n16681), .ZN(n16679) );
  OAI21_X1 U11210 ( .B1(\pipeline/immediate_to_exe [6]), .B2(n17327), .A(
        n16679), .ZN(n15538) );
  XNOR2_X1 U11208 ( .A(n17381), .B(n15537), .ZN(n16676) );
  AOI22_X1 U11206 ( .A1(n17663), .A2(\pipeline/Alu_Out_Addr_to_mem[6] ), .B1(
        n17664), .B2(n13842), .ZN(n16678) );
  NAND2_X1 U11204 ( .A1(n16676), .A2(\pipeline/stageE/input1_to_ALU [6]), .ZN(
        n15525) );
  NAND2_X1 U11203 ( .A1(n16677), .A2(\pipeline/stageE/input1_to_ALU [5]), .ZN(
        n15540) );
  AOI22_X1 U11281 ( .A1(n17663), .A2(\pipeline/Alu_Out_Addr_to_mem[7] ), .B1(
        n17664), .B2(n13839), .ZN(n16713) );
  NOR2_X1 U11286 ( .A1(\pipeline/EXE_controls_in_EXEcute [0]), .A2(n13841), 
        .ZN(n16715) );
  AOI22_X1 U11285 ( .A1(n16607), .A2(\pipeline/Alu_Out_Addr_to_mem[7] ), .B1(
        n17670), .B2(\pipeline/data_to_RF_from_WB[7] ), .ZN(n16716) );
  OAI21_X1 U11284 ( .B1(n17120), .B2(n16715), .A(n16716), .ZN(n16714) );
  OAI21_X1 U11283 ( .B1(\pipeline/immediate_to_exe [7]), .B2(n17327), .A(
        n16714), .ZN(n15512) );
  NOR2_X1 U11293 ( .A1(\pipeline/EXE_controls_in_EXEcute [0]), .A2(n13875), 
        .ZN(n16718) );
  AOI22_X1 U11292 ( .A1(n16607), .A2(\pipeline/Alu_Out_Addr_to_mem[8] ), .B1(
        n17670), .B2(\pipeline/data_to_RF_from_WB[8] ), .ZN(n16719) );
  OAI21_X1 U11291 ( .B1(n17120), .B2(n16718), .A(n16719), .ZN(n16717) );
  OAI21_X1 U11290 ( .B1(\pipeline/immediate_to_exe [8]), .B2(n17327), .A(
        n16717), .ZN(n15498) );
  XNOR2_X1 U11288 ( .A(n17381), .B(n15505), .ZN(n16672) );
  NAND2_X1 U11196 ( .A1(n16672), .A2(\pipeline/stageE/input1_to_ALU [8]), .ZN(
        n15479) );
  NOR2_X1 U11191 ( .A1(\pipeline/EXE_controls_in_EXEcute [0]), .A2(n13822), 
        .ZN(n16669) );
  AOI22_X1 U11190 ( .A1(n17665), .A2(\pipeline/Alu_Out_Addr_to_mem[9] ), .B1(
        n17123), .B2(\pipeline/data_to_RF_from_WB[9] ), .ZN(n16670) );
  OAI21_X1 U11189 ( .B1(n17120), .B2(n16669), .A(n16670), .ZN(n16668) );
  OAI21_X1 U11188 ( .B1(\pipeline/immediate_to_exe [9]), .B2(n17327), .A(
        n16668), .ZN(n15492) );
  XNOR2_X1 U11186 ( .A(n17381), .B(n15491), .ZN(n16667) );
  NOR2_X1 U11185 ( .A1(\pipeline/stageE/input1_to_ALU [9]), .A2(n16667), .ZN(
        n15477) );
  NOR2_X1 U11304 ( .A1(\pipeline/EXE_controls_in_EXEcute [0]), .A2(n13827), 
        .ZN(n16723) );
  AOI22_X1 U11303 ( .A1(n17665), .A2(\pipeline/Alu_Out_Addr_to_mem[10] ), .B1(
        n17670), .B2(\pipeline/data_to_RF_from_WB[10] ), .ZN(n16724) );
  OAI21_X1 U11302 ( .B1(n17120), .B2(n16723), .A(n16724), .ZN(n16722) );
  OAI21_X1 U11301 ( .B1(\pipeline/immediate_to_exe [10]), .B2(n17327), .A(
        n16722), .ZN(n15474) );
  AOI22_X1 U11299 ( .A1(n17663), .A2(\pipeline/Alu_Out_Addr_to_mem[10] ), .B1(
        n17664), .B2(n13826), .ZN(n16721) );
  NAND2_X1 U11181 ( .A1(n16666), .A2(\pipeline/stageE/input1_to_ALU [10]), 
        .ZN(n15463) );
  NAND2_X1 U11182 ( .A1(n16667), .A2(\pipeline/stageE/input1_to_ALU [9]), .ZN(
        n15480) );
  AOI22_X1 U11306 ( .A1(n17663), .A2(\pipeline/Alu_Out_Addr_to_mem[11] ), .B1(
        n17664), .B2(n13823), .ZN(n16725) );
  NOR2_X1 U11311 ( .A1(\pipeline/EXE_controls_in_EXEcute [0]), .A2(n13825), 
        .ZN(n16727) );
  AOI22_X1 U11310 ( .A1(n16607), .A2(\pipeline/Alu_Out_Addr_to_mem[11] ), .B1(
        n17670), .B2(\pipeline/data_to_RF_from_WB[11] ), .ZN(n16728) );
  OAI21_X1 U11309 ( .B1(n17120), .B2(n16727), .A(n16728), .ZN(n16726) );
  OAI21_X1 U11308 ( .B1(\pipeline/immediate_to_exe [11]), .B2(n17327), .A(
        n16726), .ZN(n15449) );
  NOR2_X1 U11178 ( .A1(\pipeline/EXE_controls_in_EXEcute [0]), .A2(n13815), 
        .ZN(n16662) );
  OAI21_X1 U11176 ( .B1(n17120), .B2(n16662), .A(n16663), .ZN(n16661) );
  OAI21_X1 U11175 ( .B1(\pipeline/immediate_to_exe [12]), .B2(n17327), .A(
        n16661), .ZN(n15435) );
  XNOR2_X1 U11173 ( .A(\pipeline/stageE/EXE_ALU/add_alu/sCout[0] ), .B(n15442), 
        .ZN(n16658) );
  AOI22_X1 U11171 ( .A1(n17663), .A2(\pipeline/Alu_Out_Addr_to_mem[12] ), .B1(
        n17664), .B2(n13814), .ZN(n16660) );
  NOR2_X1 U11168 ( .A1(n16658), .A2(n17080), .ZN(n15431) );
  NOR2_X1 U11165 ( .A1(\pipeline/stageE/input1_to_ALU [13]), .A2(n16659), .ZN(
        n15414) );
  NAND2_X1 U11163 ( .A1(n17080), .A2(n16658), .ZN(n15430) );
  NOR2_X1 U11162 ( .A1(\pipeline/EXE_controls_in_EXEcute [0]), .A2(n13874), 
        .ZN(n16655) );
  AOI22_X1 U11161 ( .A1(n17665), .A2(\pipeline/Alu_Out_Addr_to_mem[14] ), .B1(
        n17670), .B2(\pipeline/data_to_RF_from_WB[14] ), .ZN(n16656) );
  OAI21_X1 U11160 ( .B1(n17120), .B2(n16655), .A(n16656), .ZN(n16654) );
  OAI21_X1 U11159 ( .B1(\pipeline/immediate_to_exe [14]), .B2(n17327), .A(
        n16654), .ZN(n15411) );
  XNOR2_X1 U11157 ( .A(\pipeline/stageE/EXE_ALU/add_alu/sCout[0] ), .B(n15410), 
        .ZN(n16651) );
  AOI22_X1 U11155 ( .A1(n17663), .A2(\pipeline/Alu_Out_Addr_to_mem[14] ), .B1(
        n17664), .B2(n13960), .ZN(n16653) );
  NAND2_X1 U11152 ( .A1(n16651), .A2(n17100), .ZN(n15400) );
  NOR2_X1 U11149 ( .A1(n17100), .A2(n16651), .ZN(n15398) );
  NOR2_X1 U11147 ( .A1(\pipeline/EXE_controls_in_EXEcute [0]), .A2(n13878), 
        .ZN(n16648) );
  AOI22_X1 U11146 ( .A1(n17665), .A2(\pipeline/Alu_Out_Addr_to_mem[15] ), .B1(
        n17670), .B2(\pipeline/data_to_RF_from_WB[15] ), .ZN(n16649) );
  OAI21_X1 U11145 ( .B1(n17120), .B2(n16648), .A(n16649), .ZN(n16647) );
  OAI21_X1 U11144 ( .B1(\pipeline/immediate_to_exe [15]), .B2(n17327), .A(
        n16647), .ZN(n15386) );
  XNOR2_X1 U11143 ( .A(n17381), .B(n15386), .ZN(n15397) );
  AOI22_X1 U11140 ( .A1(n17663), .A2(\pipeline/Alu_Out_Addr_to_mem[17] ), .B1(
        n17664), .B2(n13946), .ZN(n16645) );
  NOR2_X1 U11138 ( .A1(\pipeline/EXE_controls_in_EXEcute [0]), .A2(n13879), 
        .ZN(n16643) );
  AOI22_X1 U11137 ( .A1(n17665), .A2(\pipeline/Alu_Out_Addr_to_mem[17] ), .B1(
        n17123), .B2(\pipeline/data_to_RF_from_WB[17] ), .ZN(n16644) );
  OAI21_X1 U11136 ( .B1(n17120), .B2(n16643), .A(n16644), .ZN(n16642) );
  OAI21_X1 U11135 ( .B1(\pipeline/immediate_to_exe [17]), .B2(n17327), .A(
        n16642), .ZN(n15363) );
  XNOR2_X1 U11133 ( .A(n17381), .B(n15362), .ZN(n16633) );
  NOR2_X1 U11132 ( .A1(\pipeline/stageE/input1_to_ALU [17]), .A2(n16633), .ZN(
        n16632) );
  OAI21_X1 U11128 ( .B1(n17105), .B2(n17426), .A(n16641), .ZN(
        \pipeline/stageE/input1_to_ALU [16]) );
  NOR2_X1 U11127 ( .A1(\pipeline/EXE_controls_in_EXEcute [0]), .A2(n13873), 
        .ZN(n16639) );
  OAI21_X1 U11125 ( .B1(n17120), .B2(n16639), .A(n16640), .ZN(n16638) );
  OAI21_X1 U11124 ( .B1(\pipeline/immediate_to_exe [16]), .B2(n17327), .A(
        n16638), .ZN(n15372) );
  XNOR2_X1 U11122 ( .A(n17381), .B(n15379), .ZN(n15369) );
  NOR2_X1 U11333 ( .A1(\pipeline/EXE_controls_in_EXEcute [0]), .A2(n13872), 
        .ZN(n16736) );
  AOI22_X1 U11332 ( .A1(n16607), .A2(\pipeline/Alu_Out_Addr_to_mem[18] ), .B1(
        n17670), .B2(\pipeline/data_to_RF_from_WB[18] ), .ZN(n16737) );
  OAI21_X1 U11331 ( .B1(n17120), .B2(n16736), .A(n16737), .ZN(n16735) );
  OAI21_X1 U11330 ( .B1(\pipeline/immediate_to_exe [18]), .B2(n17327), .A(
        n16735), .ZN(n15346) );
  NOR2_X1 U11115 ( .A1(\pipeline/EXE_controls_in_EXEcute [0]), .A2(n13880), 
        .ZN(n16635) );
  AOI22_X1 U11114 ( .A1(n17666), .A2(\pipeline/Alu_Out_Addr_to_mem[19] ), .B1(
        n17670), .B2(\pipeline/data_to_RF_from_WB[19] ), .ZN(n16636) );
  OAI21_X1 U11113 ( .B1(n17120), .B2(n16635), .A(n16636), .ZN(n16634) );
  OAI21_X1 U11112 ( .B1(\pipeline/immediate_to_exe [19]), .B2(n17327), .A(
        n16634), .ZN(n15331) );
  XNOR2_X1 U11110 ( .A(n17381), .B(n15330), .ZN(n15314) );
  NAND2_X1 U11100 ( .A1(n17097), .A2(n15332), .ZN(n15316) );
  NOR2_X1 U11349 ( .A1(\pipeline/EXE_controls_in_EXEcute [0]), .A2(n13881), 
        .ZN(n16744) );
  AOI22_X1 U11348 ( .A1(n17666), .A2(\pipeline/Alu_Out_Addr_to_mem[21] ), .B1(
        n17670), .B2(\pipeline/data_to_RF_from_WB[21] ), .ZN(n16745) );
  OAI21_X1 U11347 ( .B1(n17120), .B2(n16744), .A(n16745), .ZN(n16743) );
  OAI21_X1 U11346 ( .B1(\pipeline/immediate_to_exe [21]), .B2(n17327), .A(
        n16743), .ZN(n15285) );
  AOI22_X1 U11344 ( .A1(n17663), .A2(\pipeline/Alu_Out_Addr_to_mem[21] ), .B1(
        n17664), .B2(n13950), .ZN(n16742) );
  NOR2_X1 U11342 ( .A1(n16626), .A2(\pipeline/stageE/input1_to_ALU [21]), .ZN(
        n15301) );
  NOR2_X1 U11341 ( .A1(\pipeline/EXE_controls_in_EXEcute [0]), .A2(n13871), 
        .ZN(n16740) );
  AOI22_X1 U11340 ( .A1(n17666), .A2(\pipeline/Alu_Out_Addr_to_mem[20] ), .B1(
        n17670), .B2(\pipeline/data_to_RF_from_WB[20] ), .ZN(n16741) );
  OAI21_X1 U11339 ( .B1(n17120), .B2(n16740), .A(n16741), .ZN(n16739) );
  OAI21_X1 U11338 ( .B1(\pipeline/immediate_to_exe [20]), .B2(n17327), .A(
        n16739), .ZN(n15312) );
  AOI22_X1 U11336 ( .A1(n17663), .A2(\pipeline/Alu_Out_Addr_to_mem[20] ), .B1(
        n17664), .B2(n13949), .ZN(n16738) );
  NOR2_X1 U11102 ( .A1(n16629), .A2(\pipeline/stageE/input1_to_ALU [20]), .ZN(
        n15298) );
  NAND2_X1 U11108 ( .A1(n15369), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/A[16] ), .ZN(n15382) );
  NAND2_X1 U11107 ( .A1(n16633), .A2(\pipeline/stageE/input1_to_ALU [17]), 
        .ZN(n15366) );
  OAI21_X1 U11106 ( .B1(n16632), .B2(n15382), .A(n15366), .ZN(n15352) );
  OAI221_X1 U11104 ( .B1(n15352), .B2(n15348), .C1(n15352), .C2(
        \pipeline/stageE/input1_to_ALU [18]), .A(n16630), .ZN(n15319) );
  NAND2_X1 U11334 ( .A1(n16629), .A2(\pipeline/stageE/input1_to_ALU [20]), 
        .ZN(n15297) );
  NAND2_X1 U11098 ( .A1(n16626), .A2(\pipeline/stageE/input1_to_ALU [21]), 
        .ZN(n15299) );
  AOI22_X1 U11359 ( .A1(n17663), .A2(\pipeline/Alu_Out_Addr_to_mem[22] ), .B1(
        n17664), .B2(n13951), .ZN(n16749) );
  NOR2_X1 U11357 ( .A1(\pipeline/EXE_controls_in_EXEcute [0]), .A2(n13870), 
        .ZN(n16747) );
  AOI22_X1 U11356 ( .A1(n17666), .A2(\pipeline/Alu_Out_Addr_to_mem[22] ), .B1(
        n17670), .B2(\pipeline/data_to_RF_from_WB[22] ), .ZN(n16748) );
  OAI21_X1 U11355 ( .B1(n17120), .B2(n16747), .A(n16748), .ZN(n16746) );
  OAI21_X1 U11354 ( .B1(\pipeline/immediate_to_exe [22]), .B2(n17327), .A(
        n16746), .ZN(n15279) );
  XNOR2_X1 U11352 ( .A(n17381), .B(n15278), .ZN(n16624) );
  NAND2_X1 U11351 ( .A1(\pipeline/stageE/input1_to_ALU [22]), .A2(n16624), 
        .ZN(n15268) );
  NOR2_X1 U11364 ( .A1(\pipeline/EXE_controls_in_EXEcute [0]), .A2(n13882), 
        .ZN(n16751) );
  OAI21_X1 U11362 ( .B1(n17120), .B2(n16751), .A(n16752), .ZN(n16750) );
  OAI21_X1 U11361 ( .B1(\pipeline/immediate_to_exe [23]), .B2(n17327), .A(
        n16750), .ZN(n15261) );
  NOR2_X1 U11095 ( .A1(n16624), .A2(\pipeline/stageE/input1_to_ALU [22]), .ZN(
        n15265) );
  AOI22_X1 U11090 ( .A1(n17663), .A2(\pipeline/Alu_Out_Addr_to_mem[24] ), .B1(
        n17664), .B2(n13963), .ZN(n16618) );
  NOR2_X1 U11087 ( .A1(\pipeline/EXE_controls_in_EXEcute [0]), .A2(n13869), 
        .ZN(n16615) );
  AOI22_X1 U11086 ( .A1(n17666), .A2(\pipeline/Alu_Out_Addr_to_mem[24] ), .B1(
        n17670), .B2(\pipeline/data_to_RF_from_WB[24] ), .ZN(n16616) );
  OAI21_X1 U11085 ( .B1(n17120), .B2(n16615), .A(n16616), .ZN(n16614) );
  OAI21_X1 U11084 ( .B1(\pipeline/immediate_to_exe [24]), .B2(n17327), .A(
        n16614), .ZN(n15246) );
  XNOR2_X1 U11082 ( .A(n17381), .B(n15245), .ZN(n15249) );
  NAND2_X1 U11080 ( .A1(n15249), .A2(\pipeline/stageE/input1_to_ALU [24]), 
        .ZN(n15250) );
  AOI22_X1 U11369 ( .A1(n17663), .A2(\pipeline/Alu_Out_Addr_to_mem[25] ), .B1(
        n17664), .B2(n13953), .ZN(n16754) );
  NOR2_X1 U11374 ( .A1(\pipeline/EXE_controls_in_EXEcute [0]), .A2(n13883), 
        .ZN(n16756) );
  OAI21_X1 U11372 ( .B1(n17120), .B2(n16756), .A(n16757), .ZN(n16755) );
  OAI21_X1 U11371 ( .B1(\pipeline/immediate_to_exe [25]), .B2(n17327), .A(
        n16755), .ZN(n15224) );
  NOR2_X1 U11382 ( .A1(\pipeline/EXE_controls_in_EXEcute [0]), .A2(n13868), 
        .ZN(n16760) );
  AOI22_X1 U11381 ( .A1(n17666), .A2(\pipeline/Alu_Out_Addr_to_mem[26] ), .B1(
        n17123), .B2(\pipeline/data_to_RF_from_WB[26] ), .ZN(n16761) );
  OAI21_X1 U11380 ( .B1(n17120), .B2(n16760), .A(n16761), .ZN(n16759) );
  OAI21_X1 U11379 ( .B1(\pipeline/immediate_to_exe [26]), .B2(n17327), .A(
        n16759), .ZN(n15216) );
  AOI22_X1 U11377 ( .A1(n17663), .A2(\pipeline/Alu_Out_Addr_to_mem[26] ), .B1(
        n17664), .B2(n13954), .ZN(n16758) );
  NOR2_X1 U11375 ( .A1(n16612), .A2(\pipeline/stageE/input1_to_ALU [26]), .ZN(
        n15220) );
  NAND2_X1 U11077 ( .A1(n16612), .A2(\pipeline/stageE/input1_to_ALU [26]), 
        .ZN(n15221) );
  AOI22_X1 U11384 ( .A1(n17663), .A2(\pipeline/Alu_Out_Addr_to_mem[27] ), .B1(
        n17664), .B2(n13955), .ZN(n16762) );
  NOR2_X1 U11389 ( .A1(\pipeline/EXE_controls_in_EXEcute [0]), .A2(n13884), 
        .ZN(n16764) );
  AOI22_X1 U11388 ( .A1(n17665), .A2(\pipeline/Alu_Out_Addr_to_mem[27] ), .B1(
        n17670), .B2(\pipeline/data_to_RF_from_WB[27] ), .ZN(n16765) );
  OAI21_X1 U11387 ( .B1(n17120), .B2(n16764), .A(n16765), .ZN(n16763) );
  OAI21_X1 U11386 ( .B1(\pipeline/immediate_to_exe [27]), .B2(n17327), .A(
        n16763), .ZN(n15202) );
  NOR2_X1 U11397 ( .A1(\pipeline/EXE_controls_in_EXEcute [0]), .A2(n13867), 
        .ZN(n16768) );
  AOI22_X1 U11396 ( .A1(n17665), .A2(\pipeline/Alu_Out_Addr_to_mem[28] ), .B1(
        n17670), .B2(\pipeline/data_to_RF_from_WB[28] ), .ZN(n16769) );
  OAI21_X1 U11395 ( .B1(n17120), .B2(n16768), .A(n16769), .ZN(n16767) );
  OAI21_X1 U11394 ( .B1(\pipeline/immediate_to_exe [28]), .B2(n17327), .A(
        n16767), .ZN(n15182) );
  NAND2_X1 U11074 ( .A1(\pipeline/stageE/input1_to_ALU [28]), .A2(n16611), 
        .ZN(n15163) );
  NAND2_X1 U9633 ( .A1(n15166), .A2(n15163), .ZN(n15191) );
  OAI21_X1 U9670 ( .B1(n15249), .B2(n17158), .A(n15250), .ZN(n15247) );
  NOR2_X1 U9652 ( .A1(n15219), .A2(n15220), .ZN(n15217) );
  OAI21_X1 U9680 ( .B1(n15265), .B2(n15267), .A(n15268), .ZN(n15264) );
  NAND2_X1 U9679 ( .A1(n17092), .A2(n15264), .ZN(n15266) );
  OAI22_X1 U9678 ( .A1(n17092), .A2(n15264), .B1(n15265), .B2(n15266), .ZN(
        n15262) );
  NAND2_X1 U9724 ( .A1(n15319), .A2(n15335), .ZN(n15334) );
  NOR2_X1 U9691 ( .A1(n15281), .A2(n15265), .ZN(n15280) );
  XNOR2_X1 U9690 ( .A(n15267), .B(n15280), .ZN(n15024) );
  XNOR2_X1 U9661 ( .A(n15233), .B(n17115), .ZN(n15020) );
  NAND2_X1 U9702 ( .A1(n15299), .A2(n15300), .ZN(n15294) );
  NOR2_X1 U9715 ( .A1(n15314), .A2(\pipeline/stageE/input1_to_ALU [19]), .ZN(
        n15318) );
  NOR2_X1 U9714 ( .A1(n15318), .A2(n15319), .ZN(n15317) );
  AOI21_X1 U9701 ( .B1(n15296), .B2(n15297), .A(n15298), .ZN(n15295) );
  NAND2_X1 U9753 ( .A1(n15382), .A2(n15383), .ZN(n15381) );
  AOI21_X1 U9777 ( .B1(n15429), .B2(n15430), .A(n15431), .ZN(n15415) );
  OAI21_X1 U9769 ( .B1(n15414), .B2(n15415), .A(n15416), .ZN(n15399) );
  OAI21_X1 U9761 ( .B1(n15398), .B2(n15399), .A(n15400), .ZN(n15395) );
  NAND2_X1 U9778 ( .A1(n15432), .A2(n15416), .ZN(n15428) );
  NAND2_X1 U9808 ( .A1(n15463), .A2(n17587), .ZN(n15475) );
  OAI21_X1 U9796 ( .B1(n15461), .B2(n15462), .A(n15463), .ZN(n15460) );
  XNOR2_X1 U9795 ( .A(n15459), .B(n15460), .ZN(n15458) );
  XNOR2_X1 U9794 ( .A(n17082), .B(n15458), .ZN(n15040) );
  NAND2_X1 U9826 ( .A1(n15479), .A2(n15509), .ZN(n15507) );
  NAND2_X1 U9837 ( .A1(n15526), .A2(n15527), .ZN(n15524) );
  NAND2_X1 U9836 ( .A1(n15524), .A2(n15525), .ZN(n15523) );
  XNOR2_X1 U9835 ( .A(n17089), .B(n15523), .ZN(n15522) );
  XNOR2_X1 U9834 ( .A(n15521), .B(n15522), .ZN(n15037) );
  NAND2_X1 U9847 ( .A1(n15527), .A2(n15525), .ZN(n15539) );
  XNOR2_X1 U9846 ( .A(n15526), .B(n15539), .ZN(n15043) );
  NOR2_X1 U9858 ( .A1(n15555), .A2(n15542), .ZN(n15554) );
  NAND2_X1 U9866 ( .A1(n15568), .A2(n15569), .ZN(n15567) );
  AOI21_X1 U9899 ( .B1(n15058), .B2(n15053), .A(n15055), .ZN(n15592) );
  AOI21_X1 U9896 ( .B1(n15594), .B2(n15053), .A(n15055), .ZN(n15593) );
  NAND2_X1 U9513 ( .A1(\pipeline/stageE/EXE_ALU/add_alu/sCout[0] ), .A2(n15058), .ZN(n15057) );
  OAI21_X1 U9512 ( .B1(\pipeline/stageE/EXE_ALU/add_alu/sCout[0] ), .B2(n15056), .A(n15057), .ZN(n15051) );
  NAND2_X1 U9510 ( .A1(n15053), .A2(n15054), .ZN(n15052) );
  XNOR2_X1 U9509 ( .A(n15051), .B(n15052), .ZN(n14948) );
  NAND2_X1 U9818 ( .A1(n15480), .A2(n15495), .ZN(n15493) );
  NAND2_X1 U9786 ( .A1(n15430), .A2(n15446), .ZN(n15444) );
  NOR2_X1 U9768 ( .A1(n15413), .A2(n15398), .ZN(n15412) );
  NOR2_X1 U9716 ( .A1(n15320), .A2(n15298), .ZN(n15313) );
  XNOR2_X1 U9712 ( .A(n15313), .B(n15296), .ZN(n15026) );
  NOR2_X1 U11407 ( .A1(\pipeline/EXE_controls_in_EXEcute [0]), .A2(n13885), 
        .ZN(n16772) );
  OAI21_X1 U11405 ( .B1(n17120), .B2(n16772), .A(n16773), .ZN(n16771) );
  OAI21_X1 U11404 ( .B1(\pipeline/immediate_to_exe [29]), .B2(n17327), .A(
        n16771), .ZN(n15169) );
  XNOR2_X1 U11402 ( .A(n17381), .B(n15176), .ZN(n16609) );
  NAND2_X1 U9613 ( .A1(n15165), .A2(n15166), .ZN(n15146) );
  NAND2_X1 U11071 ( .A1(\pipeline/stageE/input1_to_ALU [29]), .A2(n16609), 
        .ZN(n15147) );
  OAI21_X1 U9612 ( .B1(n15163), .B2(n15164), .A(n15147), .ZN(n15162) );
  NOR2_X1 U11415 ( .A1(\pipeline/EXE_controls_in_EXEcute [0]), .A2(n13866), 
        .ZN(n16775) );
  AOI22_X1 U11414 ( .A1(n17665), .A2(\pipeline/Alu_Out_Addr_to_mem[30] ), .B1(
        n17123), .B2(\pipeline/data_to_RF_from_WB[30] ), .ZN(n16776) );
  OAI21_X1 U11413 ( .B1(n17642), .B2(n16775), .A(n16776), .ZN(n16774) );
  OAI21_X1 U11412 ( .B1(\pipeline/immediate_to_exe [30]), .B2(n17327), .A(
        n16774), .ZN(n15150) );
  XNOR2_X1 U11410 ( .A(\pipeline/stageE/EXE_ALU/add_alu/sCout[0] ), .B(n15157), 
        .ZN(n16608) );
  AOI22_X1 U11435 ( .A1(n16619), .A2(\pipeline/Alu_Out_Addr_to_mem[30] ), .B1(
        n17664), .B2(n13957), .ZN(n16792) );
  NAND2_X1 U11409 ( .A1(n17083), .A2(n16608), .ZN(n15142) );
  NAND2_X1 U9608 ( .A1(n15138), .A2(n15142), .ZN(n15160) );
  AOI22_X1 U11439 ( .A1(n17663), .A2(\pipeline/Alu_Out_Addr_to_mem[31] ), .B1(
        n17664), .B2(n13966), .ZN(n16793) );
  NOR2_X1 U11067 ( .A1(\pipeline/EXE_controls_in_EXEcute [0]), .A2(n13886), 
        .ZN(n16605) );
  AOI22_X1 U11066 ( .A1(n17666), .A2(\pipeline/Alu_Out_Addr_to_mem[31] ), .B1(
        n17670), .B2(\pipeline/data_to_RF_from_WB[31] ), .ZN(n16606) );
  OAI21_X1 U11065 ( .B1(n17642), .B2(n16605), .A(n16606), .ZN(n16603) );
  OAI21_X1 U11064 ( .B1(\pipeline/immediate_to_exe [31]), .B2(n17327), .A(
        n16603), .ZN(n15134) );
  NOR2_X1 U9882 ( .A1(n17381), .A2(n15586), .ZN(n15583) );
  NAND2_X1 U9879 ( .A1(n15583), .A2(n17405), .ZN(n15584) );
  NAND2_X1 U9881 ( .A1(\pipeline/EXE_controls_in_EXEcute [3]), .A2(n15583), 
        .ZN(n15581) );
  NAND2_X1 U9876 ( .A1(\pipeline/EXE_controls_in_EXEcute [2]), .A2(n15583), 
        .ZN(n15582) );
  NOR2_X1 U10219 ( .A1(n15834), .A2(n14127), .ZN(n15607) );
  AOI22_X1 U10053 ( .A1(\pipeline/stageF/PC_plus4/N35 ), .A2(n17108), .B1(
        n17674), .B2(n13865), .ZN(n15689) );
  AOI22_X1 U10051 ( .A1(\pipeline/stageD/target_Jump_temp [28]), .A2(n15607), 
        .B1(n17106), .B2(n15692), .ZN(n15690) );
  AOI22_X1 U10050 ( .A1(\pipeline/data_to_RF_from_WB[28] ), .A2(n17332), .B1(
        \pipeline/Alu_Out_Addr_to_mem[28] ), .B2(n17330), .ZN(n15691) );
  AOI22_X1 U10059 ( .A1(\pipeline/stageF/PC_plus4/N34 ), .A2(n17108), .B1(
        n15611), .B2(n13864), .ZN(n15694) );
  AOI22_X1 U10057 ( .A1(\pipeline/stageD/target_Jump_temp [27]), .A2(n17676), 
        .B1(n17106), .B2(n15697), .ZN(n15695) );
  AOI22_X1 U10056 ( .A1(\pipeline/data_to_RF_from_WB[27] ), .A2(n17332), .B1(
        \pipeline/Alu_Out_Addr_to_mem[27] ), .B2(n17330), .ZN(n15696) );
  NAND2_X1 U9892 ( .A1(n17421), .A2(n14995), .ZN(n15588) );
  AOI22_X1 U9596 ( .A1(n17150), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N38 ), 
        .B1(n17149), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N70 ), .ZN(n15128)
         );
  AOI22_X1 U9595 ( .A1(n17680), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N168 ), 
        .B1(n17126), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N136 ), .ZN(n15129) );
  AOI22_X1 U9594 ( .A1(n17419), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N233 ), 
        .B1(n17360), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N265 ), .ZN(n15130) );
  NAND4_X1 U9593 ( .A1(n15128), .A2(n15129), .A3(n15130), .A4(n15131), .ZN(
        n15127) );
  NAND2_X1 U9591 ( .A1(n15124), .A2(n15125), .ZN(\pipeline/EXMEM_stage/N38 )
         );
  NOR2_X1 U9607 ( .A1(\pipeline/stageE/input1_to_ALU [30]), .A2(n15150), .ZN(
        n15151) );
  AOI22_X1 U9606 ( .A1(n17150), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N37 ), 
        .B1(n17149), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N69 ), .ZN(n15154)
         );
  AOI22_X1 U9605 ( .A1(n17359), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N167 ), 
        .B1(n14964), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N135 ), .ZN(n15155) );
  AOI22_X1 U9604 ( .A1(n17419), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N232 ), 
        .B1(n17360), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N264 ), .ZN(n15156) );
  AOI211_X1 U9603 ( .C1(n14954), .C2(n15151), .A(n15152), .B(n15153), .ZN(
        n15148) );
  OAI211_X1 U9602 ( .C1(n15009), .C2(n14949), .A(n15148), .B(n15149), .ZN(
        \pipeline/EXMEM_stage/N37 ) );
  AOI22_X1 U10065 ( .A1(\pipeline/stageF/PC_plus4/N33 ), .A2(n17108), .B1(
        n17674), .B2(n13863), .ZN(n15699) );
  AOI22_X1 U10063 ( .A1(\pipeline/stageD/target_Jump_temp [26]), .A2(n17676), 
        .B1(n17106), .B2(n15702), .ZN(n15700) );
  AOI22_X1 U10062 ( .A1(\pipeline/data_to_RF_from_WB[26] ), .A2(n17332), .B1(
        \pipeline/Alu_Out_Addr_to_mem[26] ), .B2(n17330), .ZN(n15701) );
  NOR2_X1 U9620 ( .A1(\pipeline/stageE/input1_to_ALU [29]), .A2(n15169), .ZN(
        n15170) );
  NAND2_X1 U9887 ( .A1(\pipeline/EXE_controls_in_EXEcute [4]), .A2(n15573), 
        .ZN(n14967) );
  AOI22_X1 U9618 ( .A1(n17150), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N36 ), 
        .B1(n17149), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N68 ), .ZN(n15173)
         );
  AOI22_X1 U9617 ( .A1(n17359), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N166 ), 
        .B1(n17126), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N134 ), .ZN(n15174) );
  AOI22_X1 U9616 ( .A1(n17419), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N231 ), 
        .B1(n17681), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N263 ), .ZN(n15175) );
  AOI211_X1 U9615 ( .C1(n14954), .C2(n15170), .A(n15171), .B(n15172), .ZN(
        n15167) );
  OAI211_X1 U9614 ( .C1(n15010), .C2(n14949), .A(n15167), .B(n15168), .ZN(
        \pipeline/EXMEM_stage/N36 ) );
  NOR2_X1 U9631 ( .A1(\pipeline/stageE/input1_to_ALU [28]), .A2(n15182), .ZN(
        n15183) );
  AOI22_X1 U9628 ( .A1(n17150), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N35 ), 
        .B1(n17149), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N67 ), .ZN(n15186)
         );
  AOI22_X1 U9627 ( .A1(n17359), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N165 ), 
        .B1(n17126), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N133 ), .ZN(n15187) );
  AOI22_X1 U9626 ( .A1(n17419), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N230 ), 
        .B1(n17681), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N262 ), .ZN(n15188) );
  AOI211_X1 U9625 ( .C1(n14954), .C2(n15183), .A(n15184), .B(n15185), .ZN(
        n15180) );
  OAI211_X1 U9624 ( .C1(n15011), .C2(n14949), .A(n15180), .B(n15181), .ZN(
        \pipeline/EXMEM_stage/N35 ) );
  AOI22_X1 U10071 ( .A1(\pipeline/stageF/PC_plus4/N32 ), .A2(n17108), .B1(
        n17674), .B2(n13862), .ZN(n15704) );
  AOI22_X1 U10069 ( .A1(\pipeline/stageD/target_Jump_temp [25]), .A2(n17675), 
        .B1(n17106), .B2(n15707), .ZN(n15705) );
  AOI22_X1 U10068 ( .A1(\pipeline/data_to_RF_from_WB[25] ), .A2(n17332), .B1(
        \pipeline/Alu_Out_Addr_to_mem[25] ), .B2(n17330), .ZN(n15706) );
  AOI22_X1 U9639 ( .A1(n17150), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N34 ), 
        .B1(n17149), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N66 ), .ZN(n15196)
         );
  AOI22_X1 U9638 ( .A1(n17359), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N164 ), 
        .B1(n17126), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N132 ), .ZN(n15197) );
  AOI22_X1 U9637 ( .A1(n17419), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N229 ), 
        .B1(n17681), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N261 ), .ZN(n15198) );
  NAND4_X1 U9636 ( .A1(n15196), .A2(n15197), .A3(n15198), .A4(n15199), .ZN(
        n15195) );
  AOI211_X1 U9635 ( .C1(n14993), .C2(n15014), .A(n15194), .B(n15195), .ZN(
        n15193) );
  NAND2_X1 U9634 ( .A1(n15192), .A2(n15193), .ZN(\pipeline/EXMEM_stage/N34 )
         );
  AOI22_X1 U9648 ( .A1(n17150), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N33 ), 
        .B1(n17149), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N65 ), .ZN(n15210)
         );
  AOI22_X1 U9647 ( .A1(n17359), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N163 ), 
        .B1(n17126), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N131 ), .ZN(n15211) );
  AOI22_X1 U9646 ( .A1(n17419), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N228 ), 
        .B1(n17681), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N260 ), .ZN(n15212) );
  NAND4_X1 U9645 ( .A1(n15210), .A2(n15211), .A3(n15212), .A4(n15213), .ZN(
        n15209) );
  AOI211_X1 U9644 ( .C1(n14993), .C2(n15015), .A(n15208), .B(n15209), .ZN(
        n15207) );
  NAND2_X1 U9643 ( .A1(n15206), .A2(n15207), .ZN(\pipeline/EXMEM_stage/N33 )
         );
  AOI22_X1 U10077 ( .A1(\pipeline/stageF/PC_plus4/N31 ), .A2(n17108), .B1(
        n17674), .B2(n13861), .ZN(n15709) );
  AOI22_X1 U10075 ( .A1(\pipeline/stageD/target_Jump_temp [24]), .A2(n17675), 
        .B1(n17106), .B2(n15712), .ZN(n15710) );
  AOI22_X1 U10074 ( .A1(\pipeline/data_to_RF_from_WB[24] ), .A2(n15605), .B1(
        \pipeline/Alu_Out_Addr_to_mem[24] ), .B2(n17330), .ZN(n15711) );
  AOI22_X1 U9676 ( .A1(n17150), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N30 ), 
        .B1(n17149), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N62 ), .ZN(n15255)
         );
  NOR2_X1 U9880 ( .A1(\pipeline/EXE_controls_in_EXEcute [2]), .A2(n15581), 
        .ZN(n14963) );
  AOI22_X1 U9675 ( .A1(n14963), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N160 ), 
        .B1(n17126), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N128 ), .ZN(n15256) );
  NOR2_X1 U9874 ( .A1(n17405), .A2(n15581), .ZN(n14962) );
  AOI22_X1 U9674 ( .A1(n14961), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N225 ), 
        .B1(n14962), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N257 ), .ZN(n15257) );
  NAND4_X1 U9673 ( .A1(n15255), .A2(n15256), .A3(n15257), .A4(n15258), .ZN(
        n15254) );
  AOI211_X1 U9672 ( .C1(n14993), .C2(n15022), .A(n15253), .B(n15254), .ZN(
        n15252) );
  NAND2_X1 U9671 ( .A1(n15251), .A2(n15252), .ZN(\pipeline/EXMEM_stage/N30 )
         );
  NOR2_X1 U9660 ( .A1(n17159), .A2(n15224), .ZN(n15225) );
  AOI22_X1 U9658 ( .A1(n17150), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N32 ), 
        .B1(n17149), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N64 ), .ZN(n15228)
         );
  AOI22_X1 U9657 ( .A1(n17359), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N162 ), 
        .B1(n14964), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N130 ), .ZN(n15229) );
  AOI22_X1 U9656 ( .A1(n14961), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N227 ), 
        .B1(n17681), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N259 ), .ZN(n15230) );
  AOI211_X1 U9655 ( .C1(n14954), .C2(n15225), .A(n15226), .B(n15227), .ZN(
        n15222) );
  OAI211_X1 U9654 ( .C1(n15020), .C2(n14949), .A(n15222), .B(n15223), .ZN(
        \pipeline/EXMEM_stage/N32 ) );
  AOI22_X1 U9723 ( .A1(n17150), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N26 ), 
        .B1(n17149), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N58 ), .ZN(n15325)
         );
  AOI22_X1 U9722 ( .A1(n14963), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N156 ), 
        .B1(n17126), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N124 ), .ZN(n15326) );
  AOI22_X1 U9721 ( .A1(n14961), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N221 ), 
        .B1(n14962), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N253 ), .ZN(n15327) );
  NAND4_X1 U9720 ( .A1(n15325), .A2(n15326), .A3(n15327), .A4(n15328), .ZN(
        n15324) );
  AOI211_X1 U9719 ( .C1(n14993), .C2(n15023), .A(n15323), .B(n15324), .ZN(
        n15322) );
  NAND2_X1 U9718 ( .A1(n15321), .A2(n15322), .ZN(\pipeline/EXMEM_stage/N26 )
         );
  AOI22_X1 U10083 ( .A1(\pipeline/stageF/PC_plus4/N30 ), .A2(n17108), .B1(
        n17674), .B2(n13860), .ZN(n15714) );
  AOI22_X1 U10081 ( .A1(\pipeline/stageD/target_Jump_temp [23]), .A2(n15607), 
        .B1(n17106), .B2(n15717), .ZN(n15715) );
  AOI22_X1 U10080 ( .A1(\pipeline/data_to_RF_from_WB[23] ), .A2(n15605), .B1(
        \pipeline/Alu_Out_Addr_to_mem[23] ), .B2(n15606), .ZN(n15716) );
  AOI22_X1 U9709 ( .A1(n14965), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N27 ), 
        .B1(n14966), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N59 ), .ZN(n15306)
         );
  AOI22_X1 U9708 ( .A1(n14963), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N157 ), 
        .B1(n17126), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N125 ), .ZN(n15307) );
  AOI22_X1 U9707 ( .A1(n17419), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N222 ), 
        .B1(n14962), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N254 ), .ZN(n15308) );
  NAND4_X1 U9706 ( .A1(n15306), .A2(n15307), .A3(n15308), .A4(n15309), .ZN(
        n15305) );
  AOI211_X1 U9705 ( .C1(n14993), .C2(n15026), .A(n15304), .B(n15305), .ZN(
        n15303) );
  NAND2_X1 U9704 ( .A1(n15302), .A2(n15303), .ZN(\pipeline/EXMEM_stage/N27 )
         );
  NOR2_X1 U9700 ( .A1(\pipeline/stageE/input1_to_ALU [21]), .A2(n15285), .ZN(
        n15286) );
  AOI22_X1 U9697 ( .A1(n17150), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N28 ), 
        .B1(n17149), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N60 ), .ZN(n15289)
         );
  AOI22_X1 U9696 ( .A1(n14963), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N158 ), 
        .B1(n17126), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N126 ), .ZN(n15290) );
  AOI22_X1 U9695 ( .A1(n14961), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N223 ), 
        .B1(n14962), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N255 ), .ZN(n15291) );
  AOI211_X1 U9694 ( .C1(n17677), .C2(n15286), .A(n15287), .B(n15288), .ZN(
        n15283) );
  OAI211_X1 U9693 ( .C1(n15017), .C2(n14949), .A(n15283), .B(n15284), .ZN(
        \pipeline/EXMEM_stage/N28 ) );
  NOR2_X1 U9793 ( .A1(\pipeline/stageE/input1_to_ALU [11]), .A2(n15449), .ZN(
        n15450) );
  AOI22_X1 U9791 ( .A1(n17150), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N18 ), 
        .B1(n17149), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N50 ), .ZN(n15453)
         );
  AOI22_X1 U9790 ( .A1(n17680), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N148 ), 
        .B1(n17126), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N116 ), .ZN(n15454) );
  AOI22_X1 U9789 ( .A1(n17419), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N213 ), 
        .B1(n17360), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N245 ), .ZN(n15455) );
  AOI211_X1 U9788 ( .C1(n17677), .C2(n15450), .A(n15451), .B(n15452), .ZN(
        n15447) );
  OAI211_X1 U9787 ( .C1(n15040), .C2(n14949), .A(n15447), .B(n15448), .ZN(
        \pipeline/EXMEM_stage/N18 ) );
  NOR2_X1 U9784 ( .A1(\pipeline/stageE/input1_to_ALU [12]), .A2(n15435), .ZN(
        n15436) );
  AOI22_X1 U9783 ( .A1(n17150), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N19 ), 
        .B1(n17149), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N51 ), .ZN(n15439)
         );
  AOI22_X1 U9782 ( .A1(n17680), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N149 ), 
        .B1(n17126), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N117 ), .ZN(n15440) );
  AOI22_X1 U9781 ( .A1(n14961), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N214 ), 
        .B1(n17360), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N246 ), .ZN(n15441) );
  AOI211_X1 U9780 ( .C1(n17677), .C2(n15436), .A(n15437), .B(n15438), .ZN(
        n15433) );
  OAI211_X1 U9779 ( .C1(n15030), .C2(n14949), .A(n15433), .B(n15434), .ZN(
        \pipeline/EXMEM_stage/N19 ) );
  AOI22_X1 U9731 ( .A1(n17150), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N25 ), 
        .B1(n17149), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N57 ), .ZN(n15340)
         );
  AOI22_X1 U9730 ( .A1(n17680), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N155 ), 
        .B1(n17126), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N123 ), .ZN(n15341) );
  AOI22_X1 U9729 ( .A1(n14961), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N220 ), 
        .B1(n17360), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N252 ), .ZN(n15342) );
  NAND4_X1 U9728 ( .A1(n15340), .A2(n15341), .A3(n15342), .A4(n15343), .ZN(
        n15339) );
  AOI211_X1 U9727 ( .C1(n14993), .C2(n15021), .A(n15338), .B(n15339), .ZN(
        n15337) );
  NAND2_X1 U9726 ( .A1(n15336), .A2(n15337), .ZN(\pipeline/EXMEM_stage/N25 )
         );
  AOI22_X1 U9775 ( .A1(n17150), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N20 ), 
        .B1(n17149), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N52 ), .ZN(n15421)
         );
  AOI22_X1 U9774 ( .A1(n17680), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N150 ), 
        .B1(n17126), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N118 ), .ZN(n15422) );
  AOI22_X1 U9773 ( .A1(n14961), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N215 ), 
        .B1(n14962), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N247 ), .ZN(n15423) );
  NAND4_X1 U9772 ( .A1(n15421), .A2(n15422), .A3(n15423), .A4(n15424), .ZN(
        n15420) );
  AOI211_X1 U9771 ( .C1(n14993), .C2(n15033), .A(n15419), .B(n15420), .ZN(
        n15418) );
  NAND2_X1 U9770 ( .A1(n15417), .A2(n15418), .ZN(\pipeline/EXMEM_stage/N20 )
         );
  NOR2_X1 U9760 ( .A1(\pipeline/stageE/input1_to_ALU [15]), .A2(n15386), .ZN(
        n15387) );
  AOI22_X1 U9758 ( .A1(n17150), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N22 ), 
        .B1(n17149), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N54 ), .ZN(n15390)
         );
  AOI22_X1 U9757 ( .A1(n14963), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N152 ), 
        .B1(n17126), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N120 ), .ZN(n15391) );
  AOI22_X1 U9756 ( .A1(n14961), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N217 ), 
        .B1(n14962), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N249 ), .ZN(n15392) );
  AOI211_X1 U9755 ( .C1(n17677), .C2(n15387), .A(n15388), .B(n15389), .ZN(
        n15384) );
  OAI211_X1 U9754 ( .C1(n15029), .C2(n14949), .A(n15384), .B(n15385), .ZN(
        \pipeline/EXMEM_stage/N22 ) );
  AOI22_X1 U9669 ( .A1(n14965), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N31 ), 
        .B1(n17149), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N63 ), .ZN(n15240)
         );
  AOI22_X1 U9668 ( .A1(n14963), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N161 ), 
        .B1(n17126), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N129 ), .ZN(n15241) );
  AOI22_X1 U9667 ( .A1(n14961), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N226 ), 
        .B1(n17681), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N258 ), .ZN(n15242) );
  NAND4_X1 U9666 ( .A1(n15240), .A2(n15241), .A3(n15242), .A4(n15243), .ZN(
        n15239) );
  AOI211_X1 U9665 ( .C1(n14993), .C2(n15013), .A(n15238), .B(n15239), .ZN(
        n15237) );
  NAND2_X1 U9664 ( .A1(n15236), .A2(n15237), .ZN(\pipeline/EXMEM_stage/N31 )
         );
  NAND2_X1 U9868 ( .A1(\pipeline/stageE/input1_to_ALU [4]), .A2(n14952), .ZN(
        n15556) );
  AOI22_X1 U9865 ( .A1(n17150), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N11 ), 
        .B1(n17149), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N43 ), .ZN(n15560)
         );
  AOI22_X1 U9864 ( .A1(n17359), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N141 ), 
        .B1(n17126), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N109 ), .ZN(n15561) );
  AOI22_X1 U9863 ( .A1(n17419), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N206 ), 
        .B1(n17681), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N238 ), .ZN(n15562) );
  NAND4_X1 U9862 ( .A1(n15560), .A2(n15561), .A3(n15562), .A4(n15563), .ZN(
        n15559) );
  AOI211_X1 U9861 ( .C1(n14993), .C2(n15041), .A(n15558), .B(n15559), .ZN(
        n15557) );
  OAI21_X1 U9860 ( .B1(\pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .B2(
        n15556), .A(n15557), .ZN(\pipeline/EXMEM_stage/N11 ) );
  AOI22_X1 U10089 ( .A1(\pipeline/stageF/PC_plus4/N29 ), .A2(n15610), .B1(
        n17674), .B2(n13859), .ZN(n15719) );
  AOI22_X1 U10087 ( .A1(\pipeline/stageD/target_Jump_temp [22]), .A2(n17676), 
        .B1(n17106), .B2(n15722), .ZN(n15720) );
  AOI22_X1 U10086 ( .A1(\pipeline/data_to_RF_from_WB[22] ), .A2(n15605), .B1(
        \pipeline/Alu_Out_Addr_to_mem[22] ), .B2(n15606), .ZN(n15721) );
  AOI22_X1 U9854 ( .A1(n17150), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N12 ), 
        .B1(n17149), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N44 ), .ZN(n15547)
         );
  AOI22_X1 U9853 ( .A1(n17359), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N142 ), 
        .B1(n17126), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N110 ), .ZN(n15548) );
  AOI22_X1 U9852 ( .A1(n17419), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N207 ), 
        .B1(n17681), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N239 ), .ZN(n15549) );
  NAND4_X1 U9851 ( .A1(n15547), .A2(n15548), .A3(n15549), .A4(n15550), .ZN(
        n15546) );
  AOI211_X1 U9850 ( .C1(n14993), .C2(n15042), .A(n15545), .B(n15546), .ZN(
        n15544) );
  NAND2_X1 U9849 ( .A1(n15543), .A2(n15544), .ZN(\pipeline/EXMEM_stage/N12 )
         );
  AOI22_X1 U9844 ( .A1(n14965), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N13 ), 
        .B1(n17149), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N45 ), .ZN(n15532)
         );
  AOI22_X1 U9843 ( .A1(n17359), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N143 ), 
        .B1(n17126), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N111 ), .ZN(n15533) );
  AOI22_X1 U9842 ( .A1(n17419), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N208 ), 
        .B1(n17681), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N240 ), .ZN(n15534) );
  NAND4_X1 U9841 ( .A1(n15532), .A2(n15533), .A3(n15534), .A4(n15535), .ZN(
        n15531) );
  AOI211_X1 U9840 ( .C1(n14993), .C2(n15043), .A(n15530), .B(n15531), .ZN(
        n15529) );
  NAND2_X1 U9839 ( .A1(n15528), .A2(n15529), .ZN(\pipeline/EXMEM_stage/N13 )
         );
  NOR2_X1 U9465 ( .A1(n12649), .A2(n17740), .ZN(n14955) );
  AOI22_X1 U9463 ( .A1(n17150), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N9 ), 
        .B1(n17149), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N41 ), .ZN(n14958)
         );
  AOI22_X1 U9462 ( .A1(n17680), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N139 ), 
        .B1(n17126), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N107 ), .ZN(n14959) );
  AOI22_X1 U9461 ( .A1(n17419), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N204 ), 
        .B1(n17360), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N236 ), .ZN(n14960) );
  AOI211_X1 U9460 ( .C1(n14954), .C2(n14955), .A(n14956), .B(n14957), .ZN(
        n14950) );
  OAI211_X1 U9459 ( .C1(n14948), .C2(n14949), .A(n14950), .B(n14951), .ZN(
        \pipeline/EXMEM_stage/N9 ) );
  NOR2_X1 U9890 ( .A1(n17739), .A2(\pipeline/stageE/input1_to_ALU [3]), .ZN(
        n15574) );
  AOI22_X1 U9883 ( .A1(n17150), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N10 ), 
        .B1(n14966), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N42 ), .ZN(n15577)
         );
  AOI22_X1 U9877 ( .A1(n17359), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N140 ), 
        .B1(n14964), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N108 ), .ZN(n15578) );
  AOI22_X1 U9873 ( .A1(n17419), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N205 ), 
        .B1(n17681), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N237 ), .ZN(n15579) );
  AOI211_X1 U9872 ( .C1(n17677), .C2(n15574), .A(n15575), .B(n15576), .ZN(
        n15570) );
  OAI211_X1 U9869 ( .C1(n15045), .C2(n14949), .A(n15570), .B(n15571), .ZN(
        \pipeline/EXMEM_stage/N10 ) );
  AOI22_X1 U9688 ( .A1(n17150), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N29 ), 
        .B1(n17149), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N61 ), .ZN(n15273)
         );
  AOI22_X1 U9687 ( .A1(n14963), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N159 ), 
        .B1(n17126), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N127 ), .ZN(n15274) );
  AOI22_X1 U9686 ( .A1(n14961), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N224 ), 
        .B1(n14962), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N256 ), .ZN(n15275) );
  NAND4_X1 U9685 ( .A1(n15273), .A2(n15274), .A3(n15275), .A4(n15276), .ZN(
        n15272) );
  AOI211_X1 U9684 ( .C1(n14993), .C2(n15024), .A(n15271), .B(n15272), .ZN(
        n15270) );
  NAND2_X1 U9683 ( .A1(n15269), .A2(n15270), .ZN(\pipeline/EXMEM_stage/N29 )
         );
  AOI22_X1 U9470 ( .A1(n17150), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N8 ), 
        .B1(n17149), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N40 ), .ZN(n14977)
         );
  AOI22_X1 U9469 ( .A1(n17680), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N138 ), 
        .B1(n17126), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N106 ), .ZN(n14978) );
  AOI22_X1 U9468 ( .A1(n17419), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N203 ), 
        .B1(n17360), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N235 ), .ZN(n14979) );
  NOR3_X1 U9467 ( .A1(n14974), .A2(n14975), .A3(n14976), .ZN(n14971) );
  OAI211_X1 U9466 ( .C1(n14970), .C2(n14949), .A(n14971), .B(n14972), .ZN(
        \pipeline/EXMEM_stage/N8 ) );
  AOI22_X1 U9742 ( .A1(n17150), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N24 ), 
        .B1(n17149), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N56 ), .ZN(n15357)
         );
  AOI22_X1 U9741 ( .A1(n17680), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N154 ), 
        .B1(n17126), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N122 ), .ZN(n15358) );
  AOI22_X1 U9740 ( .A1(n14961), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N219 ), 
        .B1(n17360), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N251 ), .ZN(n15359) );
  NAND4_X1 U9739 ( .A1(n15357), .A2(n15358), .A3(n15359), .A4(n15360), .ZN(
        n15356) );
  AOI211_X1 U9738 ( .C1(n14993), .C2(n15025), .A(n15355), .B(n15356), .ZN(
        n15354) );
  NAND2_X1 U9737 ( .A1(n15353), .A2(n15354), .ZN(\pipeline/EXMEM_stage/N24 )
         );
  NOR2_X1 U9752 ( .A1(\pipeline/stageE/EXE_ALU/alu_shift/C48/A[16] ), .A2(
        n15372), .ZN(n15373) );
  AOI22_X1 U9750 ( .A1(n17150), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N23 ), 
        .B1(n14966), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N55 ), .ZN(n15376)
         );
  AOI22_X1 U9749 ( .A1(n14963), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N153 ), 
        .B1(n14964), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N121 ), .ZN(n15377) );
  AOI22_X1 U9748 ( .A1(n14961), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N218 ), 
        .B1(n17681), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N250 ), .ZN(n15378) );
  AOI211_X1 U9747 ( .C1(n17677), .C2(n15373), .A(n15374), .B(n15375), .ZN(
        n15370) );
  OAI211_X1 U9746 ( .C1(n15032), .C2(n14949), .A(n15370), .B(n15371), .ZN(
        \pipeline/EXMEM_stage/N23 ) );
  NOR2_X1 U9825 ( .A1(\pipeline/stageE/input1_to_ALU [8]), .A2(n15498), .ZN(
        n15499) );
  AOI22_X1 U9823 ( .A1(n17150), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N15 ), 
        .B1(n17149), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N47 ), .ZN(n15502)
         );
  AOI22_X1 U9822 ( .A1(n17359), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N145 ), 
        .B1(n17126), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N113 ), .ZN(n15503) );
  AOI22_X1 U9821 ( .A1(n17419), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N210 ), 
        .B1(n17360), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N242 ), .ZN(n15504) );
  AOI211_X1 U9820 ( .C1(n17677), .C2(n15499), .A(n15500), .B(n15501), .ZN(
        n15496) );
  OAI211_X1 U9819 ( .C1(n15039), .C2(n14949), .A(n15496), .B(n15497), .ZN(
        \pipeline/EXMEM_stage/N15 ) );
  AOI22_X1 U9803 ( .A1(n17150), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N17 ), 
        .B1(n17149), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N49 ), .ZN(n15468)
         );
  AOI22_X1 U9802 ( .A1(n17680), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N147 ), 
        .B1(n17126), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N115 ), .ZN(n15469) );
  AOI22_X1 U9801 ( .A1(n17419), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N212 ), 
        .B1(n17360), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N244 ), .ZN(n15470) );
  NAND4_X1 U9800 ( .A1(n15468), .A2(n15469), .A3(n15470), .A4(n15471), .ZN(
        n15467) );
  AOI211_X1 U9799 ( .C1(n14993), .C2(n15034), .A(n15466), .B(n15467), .ZN(
        n15465) );
  NAND2_X1 U9798 ( .A1(n15464), .A2(n15465), .ZN(\pipeline/EXMEM_stage/N17 )
         );
  AOI22_X1 U9815 ( .A1(n17150), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N16 ), 
        .B1(n17149), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N48 ), .ZN(n15486)
         );
  AOI22_X1 U9814 ( .A1(n17680), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N146 ), 
        .B1(n17126), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N114 ), .ZN(n15487) );
  AOI22_X1 U9813 ( .A1(n17419), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N211 ), 
        .B1(n17360), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N243 ), .ZN(n15488) );
  NAND4_X1 U9812 ( .A1(n15486), .A2(n15487), .A3(n15488), .A4(n15489), .ZN(
        n15485) );
  AOI211_X1 U9811 ( .C1(n14993), .C2(n15035), .A(n15484), .B(n15485), .ZN(
        n15483) );
  NAND2_X1 U9810 ( .A1(n15482), .A2(n15483), .ZN(\pipeline/EXMEM_stage/N16 )
         );
  NOR2_X1 U9833 ( .A1(\pipeline/stageE/input1_to_ALU [7]), .A2(n15512), .ZN(
        n15513) );
  AOI22_X1 U9831 ( .A1(n17150), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N14 ), 
        .B1(n17149), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N46 ), .ZN(n15516)
         );
  AOI22_X1 U9830 ( .A1(n17359), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N144 ), 
        .B1(n14964), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N112 ), .ZN(n15517) );
  AOI22_X1 U9829 ( .A1(n17419), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N209 ), 
        .B1(n17360), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N241 ), .ZN(n15518) );
  AOI211_X1 U9828 ( .C1(n17677), .C2(n15513), .A(n15514), .B(n15515), .ZN(
        n15510) );
  OAI211_X1 U9827 ( .C1(n15037), .C2(n14949), .A(n15510), .B(n15511), .ZN(
        \pipeline/EXMEM_stage/N14 ) );
  AOI22_X1 U9767 ( .A1(n17150), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N21 ), 
        .B1(n17149), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N53 ), .ZN(n15405)
         );
  AOI22_X1 U9766 ( .A1(n17680), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N151 ), 
        .B1(n17126), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N119 ), .ZN(n15406) );
  AOI22_X1 U9765 ( .A1(n14961), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N216 ), 
        .B1(n14962), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N248 ), .ZN(n15407) );
  NAND4_X1 U9764 ( .A1(n15405), .A2(n15406), .A3(n15407), .A4(n15408), .ZN(
        n15404) );
  AOI211_X1 U9763 ( .C1(n14993), .C2(n15027), .A(n15403), .B(n15404), .ZN(
        n15402) );
  NAND2_X1 U9762 ( .A1(n15401), .A2(n15402), .ZN(\pipeline/EXMEM_stage/N21 )
         );
  AOI22_X1 U10095 ( .A1(\pipeline/stageF/PC_plus4/N28 ), .A2(n15610), .B1(
        n17674), .B2(n13858), .ZN(n15724) );
  AOI22_X1 U10093 ( .A1(\pipeline/stageD/target_Jump_temp [21]), .A2(n17675), 
        .B1(n15608), .B2(n15727), .ZN(n15725) );
  AOI22_X1 U10092 ( .A1(\pipeline/data_to_RF_from_WB[21] ), .A2(n15605), .B1(
        \pipeline/Alu_Out_Addr_to_mem[21] ), .B2(n15606), .ZN(n15726) );
  AOI22_X1 U9981 ( .A1(\pipeline/inst_IFID_DEC[31] ), .A2(n15600), .B1(n17673), 
        .B2(InstrFetched[31]), .ZN(n15653) );
  AOI22_X1 U9973 ( .A1(\pipeline/inst_IFID_DEC[27] ), .A2(n15600), .B1(n17107), 
        .B2(InstrFetched[27]), .ZN(n15649) );
  AOI22_X1 U9969 ( .A1(\pipeline/stageD/offset_jump_sign_ext [31]), .A2(n15600), .B1(n17107), .B2(InstrFetched[25]), .ZN(n15645) );
  AOI22_X1 U9961 ( .A1(\pipeline/stageD/offset_jump_sign_ext [21]), .A2(n17671), .B1(n17107), .B2(InstrFetched[21]), .ZN(n15641) );
  AOI22_X1 U9977 ( .A1(\pipeline/inst_IFID_DEC[29] ), .A2(n15600), .B1(n17673), 
        .B2(InstrFetched[29]), .ZN(n15651) );
  AOI22_X1 U9963 ( .A1(\pipeline/stageD/offset_jump_sign_ext [22]), .A2(n15600), .B1(n17107), .B2(InstrFetched[22]), .ZN(n15642) );
  AOI22_X1 U10145 ( .A1(n15600), .A2(\pipeline/nextPC_IFID_DEC[8] ), .B1(
        n17673), .B2(\pipeline/stageF/PC_plus4/N15 ), .ZN(n15768) );
  AOI22_X1 U10156 ( .A1(n15600), .A2(\pipeline/nextPC_IFID_DEC[3] ), .B1(
        n17673), .B2(\pipeline/stageF/PC_plus4/N10 ), .ZN(n15778) );
  AOI22_X1 U10067 ( .A1(n15600), .A2(\pipeline/nextPC_IFID_DEC[26] ), .B1(
        n17673), .B2(\pipeline/stageF/PC_plus4/N33 ), .ZN(n15703) );
  AOI22_X1 U9941 ( .A1(n15600), .A2(\pipeline/stageD/offset_to_jump_temp [10]), 
        .B1(n17673), .B2(InstrFetched[10]), .ZN(n15631) );
  AOI22_X1 U9965 ( .A1(\pipeline/stageD/offset_jump_sign_ext [23]), .A2(n17671), .B1(n17107), .B2(InstrFetched[23]), .ZN(n15643) );
  AOI22_X1 U10055 ( .A1(n15600), .A2(\pipeline/nextPC_IFID_DEC[28] ), .B1(
        n15601), .B2(\pipeline/stageF/PC_plus4/N35 ), .ZN(n15693) );
  AOI22_X1 U10198 ( .A1(n17671), .A2(\pipeline/nextPC_IFID_DEC[10] ), .B1(
        n17107), .B2(\pipeline/stageF/PC_plus4/N17 ), .ZN(n15813) );
  AOI22_X1 U10174 ( .A1(n15600), .A2(\pipeline/nextPC_IFID_DEC[5] ), .B1(
        n15601), .B2(\pipeline/stageF/PC_plus4/N12 ), .ZN(n15793) );
  AOI22_X1 U9931 ( .A1(n17671), .A2(\pipeline/stageD/offset_to_jump_temp [5]), 
        .B1(n17107), .B2(InstrFetched[5]), .ZN(n15626) );
  AOI22_X1 U10091 ( .A1(n15600), .A2(\pipeline/nextPC_IFID_DEC[22] ), .B1(
        n17107), .B2(\pipeline/stageF/PC_plus4/N29 ), .ZN(n15723) );
  AOI22_X1 U10109 ( .A1(n15600), .A2(\pipeline/nextPC_IFID_DEC[19] ), .B1(
        n17107), .B2(\pipeline/stageF/PC_plus4/N26 ), .ZN(n15738) );
  AOI22_X1 U9953 ( .A1(n15600), .A2(\pipeline/stageD/offset_jump_sign_ext [17]), .B1(n15601), .B2(InstrFetched[17]), .ZN(n15637) );
  AOI22_X1 U10168 ( .A1(n15600), .A2(\pipeline/nextPC_IFID_DEC[4] ), .B1(
        n15601), .B2(\pipeline/stageF/PC_plus4/N11 ), .ZN(n15788) );
  AOI22_X1 U9929 ( .A1(n17671), .A2(\pipeline/stageD/offset_to_jump_temp [4]), 
        .B1(n17107), .B2(InstrFetched[4]), .ZN(n15625) );
  AOI22_X1 U10079 ( .A1(n17671), .A2(\pipeline/nextPC_IFID_DEC[24] ), .B1(
        n17673), .B2(\pipeline/stageF/PC_plus4/N31 ), .ZN(n15713) );
  AOI22_X1 U10139 ( .A1(n17671), .A2(\pipeline/nextPC_IFID_DEC[13] ), .B1(
        n17673), .B2(\pipeline/stageF/PC_plus4/N20 ), .ZN(n15763) );
  AOI22_X1 U9905 ( .A1(n17671), .A2(\pipeline/stageD/offset_to_jump_temp [14]), 
        .B1(n17673), .B2(InstrFetched[14]), .ZN(n15599) );
  AOI22_X1 U9951 ( .A1(n17671), .A2(\pipeline/stageD/offset_jump_sign_ext [16]), .B1(n17673), .B2(InstrFetched[16]), .ZN(n15636) );
  AOI22_X1 U10162 ( .A1(n17671), .A2(\pipeline/nextPC_IFID_DEC[7] ), .B1(
        n17673), .B2(\pipeline/stageF/PC_plus4/N14 ), .ZN(n15783) );
  AOI22_X1 U10230 ( .A1(n17671), .A2(\pipeline/nextPC_IFID_DEC[30] ), .B1(
        n17107), .B2(\pipeline/stageF/PC_plus4/N37 ), .ZN(n15837) );
  AOI22_X1 U9957 ( .A1(n17671), .A2(\pipeline/stageD/offset_jump_sign_ext [19]), .B1(n17107), .B2(InstrFetched[19]), .ZN(n15639) );
  AOI22_X1 U10210 ( .A1(n17671), .A2(\pipeline/nextPC_IFID_DEC[2] ), .B1(
        n17107), .B2(\pipeline/stageF/PC_plus4/N9 ), .ZN(n15823) );
  AOI22_X1 U9959 ( .A1(n17671), .A2(\pipeline/stageD/offset_jump_sign_ext [20]), .B1(n17107), .B2(InstrFetched[20]), .ZN(n15640) );
  AOI22_X1 U10127 ( .A1(n17671), .A2(\pipeline/nextPC_IFID_DEC[15] ), .B1(
        n17107), .B2(\pipeline/stageF/PC_plus4/N22 ), .ZN(n15753) );
  AOI22_X1 U10121 ( .A1(n17671), .A2(\pipeline/nextPC_IFID_DEC[17] ), .B1(
        n17672), .B2(\pipeline/stageF/PC_plus4/N24 ), .ZN(n15748) );
  AOI22_X1 U10103 ( .A1(n17671), .A2(\pipeline/nextPC_IFID_DEC[20] ), .B1(
        n17107), .B2(\pipeline/stageF/PC_plus4/N27 ), .ZN(n15733) );
  AOI22_X1 U9939 ( .A1(n17671), .A2(\pipeline/stageD/offset_to_jump_temp [9]), 
        .B1(n17107), .B2(InstrFetched[9]), .ZN(n15630) );
  AOI22_X1 U9947 ( .A1(n15600), .A2(\pipeline/stageD/offset_to_jump_temp [13]), 
        .B1(n17673), .B2(InstrFetched[13]), .ZN(n15634) );
  AOI22_X1 U9943 ( .A1(n15600), .A2(\pipeline/stageD/offset_to_jump_temp [11]), 
        .B1(n17673), .B2(InstrFetched[11]), .ZN(n15632) );
  AOI22_X1 U10073 ( .A1(n15600), .A2(\pipeline/nextPC_IFID_DEC[25] ), .B1(
        n17673), .B2(\pipeline/stageF/PC_plus4/N32 ), .ZN(n15708) );
  AOI22_X1 U10097 ( .A1(n15600), .A2(\pipeline/nextPC_IFID_DEC[21] ), .B1(
        n17672), .B2(\pipeline/stageF/PC_plus4/N28 ), .ZN(n15728) );
  AOI22_X1 U9923 ( .A1(n17671), .A2(\pipeline/stageD/offset_to_jump_temp [1]), 
        .B1(n15601), .B2(InstrFetched[1]), .ZN(n15622) );
  AOI22_X1 U9933 ( .A1(n17671), .A2(\pipeline/stageD/offset_to_jump_temp [6]), 
        .B1(n17107), .B2(InstrFetched[6]), .ZN(n15627) );
  AOI22_X1 U9945 ( .A1(n15600), .A2(\pipeline/stageD/offset_to_jump_temp [12]), 
        .B1(n15601), .B2(InstrFetched[12]), .ZN(n15633) );
  AOI22_X1 U10061 ( .A1(n15600), .A2(\pipeline/nextPC_IFID_DEC[27] ), .B1(
        n15601), .B2(\pipeline/stageF/PC_plus4/N34 ), .ZN(n15698) );
  AOI22_X1 U10204 ( .A1(n17671), .A2(\pipeline/nextPC_IFID_DEC[12] ), .B1(
        n17107), .B2(\pipeline/stageF/PC_plus4/N19 ), .ZN(n15818) );
  AOI22_X1 U10192 ( .A1(n17671), .A2(\pipeline/nextPC_IFID_DEC[9] ), .B1(
        n17672), .B2(\pipeline/stageF/PC_plus4/N16 ), .ZN(n15808) );
  AOI22_X1 U10186 ( .A1(n15600), .A2(\pipeline/nextPC_IFID_DEC[11] ), .B1(
        n17107), .B2(\pipeline/stageF/PC_plus4/N18 ), .ZN(n15803) );
  AOI22_X1 U10226 ( .A1(n15600), .A2(\pipeline/nextPC_IFID_DEC[1] ), .B1(
        n17107), .B2(\pipeline/stageF/PC_plus4/N8 ), .ZN(n15835) );
  AOI22_X1 U9955 ( .A1(n15600), .A2(\pipeline/stageD/offset_jump_sign_ext [18]), .B1(n17673), .B2(InstrFetched[18]), .ZN(n15638) );
  AOI22_X1 U9949 ( .A1(n15600), .A2(\pipeline/stageD/offset_to_jump_temp [15]), 
        .B1(n17673), .B2(InstrFetched[15]), .ZN(n15635) );
  AOI22_X1 U10101 ( .A1(\pipeline/stageF/PC_plus4/N27 ), .A2(n15610), .B1(
        n17674), .B2(n13857), .ZN(n15729) );
  AOI22_X1 U10099 ( .A1(\pipeline/stageD/target_Jump_temp [20]), .A2(n15607), 
        .B1(n17106), .B2(n15732), .ZN(n15730) );
  AOI22_X1 U10098 ( .A1(\pipeline/data_to_RF_from_WB[20] ), .A2(n15605), .B1(
        \pipeline/Alu_Out_Addr_to_mem[20] ), .B2(n15606), .ZN(n15731) );
  AOI22_X1 U10202 ( .A1(\pipeline/stageF/PC_plus4/N19 ), .A2(n17108), .B1(
        n17674), .B2(n13813), .ZN(n15814) );
  AOI22_X1 U10200 ( .A1(\pipeline/stageD/target_Jump_temp [12]), .A2(n17675), 
        .B1(n17106), .B2(n15817), .ZN(n15815) );
  AOI22_X1 U10199 ( .A1(\pipeline/data_to_RF_from_WB[12] ), .A2(n17332), .B1(
        \pipeline/Alu_Out_Addr_to_mem[12] ), .B2(n17330), .ZN(n15816) );
  AOI22_X1 U10143 ( .A1(\pipeline/stageF/PC_plus4/N15 ), .A2(n17108), .B1(
        n17674), .B2(n13850), .ZN(n15764) );
  AOI22_X1 U10141 ( .A1(\pipeline/stageD/target_Jump_temp [8]), .A2(n17676), 
        .B1(n17106), .B2(n15767), .ZN(n15765) );
  AOI22_X1 U10140 ( .A1(\pipeline/data_to_RF_from_WB[8] ), .A2(n17333), .B1(
        \pipeline/Alu_Out_Addr_to_mem[8] ), .B2(n15606), .ZN(n15766) );
  AOI22_X1 U10113 ( .A1(\pipeline/stageF/PC_plus4/N25 ), .A2(n17108), .B1(
        n17674), .B2(n13855), .ZN(n15739) );
  AOI22_X1 U10111 ( .A1(\pipeline/stageD/target_Jump_temp [18]), .A2(n17675), 
        .B1(n17106), .B2(n15742), .ZN(n15740) );
  AOI22_X1 U10110 ( .A1(\pipeline/data_to_RF_from_WB[18] ), .A2(n15605), .B1(
        \pipeline/Alu_Out_Addr_to_mem[18] ), .B2(n15606), .ZN(n15741) );
  AOI22_X1 U10125 ( .A1(\pipeline/stageF/PC_plus4/N22 ), .A2(n17108), .B1(
        n15611), .B2(n13853), .ZN(n15749) );
  AOI22_X1 U10123 ( .A1(\pipeline/stageD/target_Jump_temp [15]), .A2(n17676), 
        .B1(n17106), .B2(n15752), .ZN(n15750) );
  AOI22_X1 U10122 ( .A1(\pipeline/data_to_RF_from_WB[15] ), .A2(n17333), .B1(
        \pipeline/Alu_Out_Addr_to_mem[15] ), .B2(n17331), .ZN(n15751) );
  AOI22_X1 U10154 ( .A1(\pipeline/stageF/PC_plus4/N10 ), .A2(n17108), .B1(
        n15611), .B2(n13845), .ZN(n15774) );
  AOI22_X1 U10152 ( .A1(\pipeline/stageD/target_Jump_temp [3]), .A2(n15607), 
        .B1(n17106), .B2(n15777), .ZN(n15775) );
  AOI22_X1 U10151 ( .A1(\pipeline/Alu_Out_Addr_to_mem[3] ), .A2(n17330), .B1(
        \pipeline/data_to_RF_from_WB[3] ), .B2(n17333), .ZN(n15776) );
  AOI22_X1 U9909 ( .A1(\pipeline/stageF/PC_plus4/N23 ), .A2(n17108), .B1(
        n17674), .B2(n13945), .ZN(n15602) );
  AOI22_X1 U9907 ( .A1(\pipeline/stageD/target_Jump_temp [16]), .A2(n17676), 
        .B1(n17106), .B2(n15609), .ZN(n15603) );
  AOI22_X1 U9906 ( .A1(\pipeline/data_to_RF_from_WB[16] ), .A2(n17333), .B1(
        \pipeline/Alu_Out_Addr_to_mem[16] ), .B2(n17331), .ZN(n15604) );
  AOI22_X1 U10196 ( .A1(\pipeline/stageF/PC_plus4/N17 ), .A2(n15610), .B1(
        n17674), .B2(n13817), .ZN(n15809) );
  AOI22_X1 U10194 ( .A1(\pipeline/stageD/target_Jump_temp [10]), .A2(n17676), 
        .B1(n17106), .B2(n15812), .ZN(n15810) );
  AOI22_X1 U10193 ( .A1(\pipeline/data_to_RF_from_WB[10] ), .A2(n17332), .B1(
        \pipeline/Alu_Out_Addr_to_mem[10] ), .B2(n17330), .ZN(n15811) );
  AOI22_X1 U10166 ( .A1(\pipeline/stageF/PC_plus4/N11 ), .A2(n17108), .B1(
        n15611), .B2(n13837), .ZN(n15784) );
  AOI22_X1 U10164 ( .A1(\pipeline/stageD/target_Jump_temp [4]), .A2(n17675), 
        .B1(n17106), .B2(n15787), .ZN(n15785) );
  AOI22_X1 U10163 ( .A1(\pipeline/data_to_RF_from_WB[4] ), .A2(n17333), .B1(
        \pipeline/Alu_Out_Addr_to_mem[4] ), .B2(n17331), .ZN(n15786) );
  AOI22_X1 U10208 ( .A1(\pipeline/stageF/PC_plus4/N9 ), .A2(n17108), .B1(
        n15611), .B2(n13810), .ZN(n15819) );
  AOI22_X1 U10206 ( .A1(\pipeline/stageD/target_Jump_temp [2]), .A2(n15607), 
        .B1(n17106), .B2(n15822), .ZN(n15820) );
  AOI22_X1 U10205 ( .A1(\pipeline/data_to_RF_from_WB[2] ), .A2(n17332), .B1(
        \pipeline/Alu_Out_Addr_to_mem[2] ), .B2(n17330), .ZN(n15821) );
  AOI22_X1 U10133 ( .A1(n15600), .A2(\pipeline/nextPC_IFID_DEC[14] ), .B1(
        n17107), .B2(\pipeline/stageF/PC_plus4/N21 ), .ZN(n15758) );
  AOI22_X1 U10115 ( .A1(n15600), .A2(\pipeline/nextPC_IFID_DEC[18] ), .B1(
        n17107), .B2(\pipeline/stageF/PC_plus4/N25 ), .ZN(n15743) );
  AOI22_X1 U9937 ( .A1(n15600), .A2(\pipeline/stageD/offset_to_jump_temp [8]), 
        .B1(n17107), .B2(InstrFetched[8]), .ZN(n15629) );
  AOI22_X1 U10228 ( .A1(n15600), .A2(\pipeline/nextPC_IFID_DEC[29] ), .B1(
        n17107), .B2(\pipeline/stageF/PC_plus4/N36 ), .ZN(n15836) );
  AOI222_X1 U10048 ( .A1(n17331), .A2(\pipeline/Alu_Out_Addr_to_mem[31] ), 
        .B1(\pipeline/stageD/target_Jump_temp [31]), .B2(n17675), .C1(n17106), 
        .C2(n15688), .ZN(n15686) );
  AOI22_X1 U10047 ( .A1(\pipeline/data_to_RF_from_WB[31] ), .A2(n17332), .B1(
        n17674), .B2(n13938), .ZN(n15687) );
  NAND2_X1 U10046 ( .A1(n15686), .A2(n15687), .ZN(n3924) );
  AOI22_X1 U10178 ( .A1(\pipeline/stageF/PC_plus4/N13 ), .A2(n17108), .B1(
        n15611), .B2(n13829), .ZN(n15794) );
  AOI22_X1 U10176 ( .A1(\pipeline/stageD/target_Jump_temp [6]), .A2(n17676), 
        .B1(n17106), .B2(n15797), .ZN(n15795) );
  AOI22_X1 U10175 ( .A1(\pipeline/data_to_RF_from_WB[6] ), .A2(n17333), .B1(
        \pipeline/Alu_Out_Addr_to_mem[6] ), .B2(n17331), .ZN(n15796) );
  AOI22_X1 U10137 ( .A1(\pipeline/stageF/PC_plus4/N20 ), .A2(n17108), .B1(
        n17674), .B2(n13851), .ZN(n15759) );
  AOI22_X1 U10135 ( .A1(\pipeline/stageD/target_Jump_temp [13]), .A2(n15607), 
        .B1(n17106), .B2(n15762), .ZN(n15760) );
  AOI22_X1 U10134 ( .A1(\pipeline/data_to_RF_from_WB[13] ), .A2(n15605), .B1(
        \pipeline/Alu_Out_Addr_to_mem[13] ), .B2(n17330), .ZN(n15761) );
  AOI22_X1 U10107 ( .A1(\pipeline/stageF/PC_plus4/N26 ), .A2(n17108), .B1(
        n17674), .B2(n13856), .ZN(n15734) );
  AOI22_X1 U10105 ( .A1(\pipeline/stageD/target_Jump_temp [19]), .A2(n17676), 
        .B1(n17106), .B2(n15737), .ZN(n15735) );
  AOI22_X1 U10104 ( .A1(\pipeline/data_to_RF_from_WB[19] ), .A2(n17333), .B1(
        \pipeline/Alu_Out_Addr_to_mem[19] ), .B2(n17331), .ZN(n15736) );
  AOI22_X1 U10148 ( .A1(\pipeline/stageF/PC_plus4/N7 ), .A2(n17108), .B1(
        n17674), .B2(n13849), .ZN(n15769) );
  AOI22_X1 U10147 ( .A1(\pipeline/stageD/target_Jump_temp [0]), .A2(n17675), 
        .B1(n17106), .B2(n15772), .ZN(n15770) );
  AOI22_X1 U10146 ( .A1(\pipeline/data_to_RF_from_WB[0] ), .A2(n17333), .B1(
        \pipeline/Alu_Out_Addr_to_mem[0] ), .B2(n15606), .ZN(n15771) );
  AOI22_X1 U10172 ( .A1(\pipeline/stageF/PC_plus4/N12 ), .A2(n17108), .B1(
        n17674), .B2(n13833), .ZN(n15789) );
  AOI22_X1 U10170 ( .A1(\pipeline/stageD/target_Jump_temp [5]), .A2(n15607), 
        .B1(n17106), .B2(n15792), .ZN(n15790) );
  AOI22_X1 U10169 ( .A1(\pipeline/data_to_RF_from_WB[5] ), .A2(n17333), .B1(
        \pipeline/Alu_Out_Addr_to_mem[5] ), .B2(n17331), .ZN(n15791) );
  AOI22_X1 U10160 ( .A1(\pipeline/stageF/PC_plus4/N14 ), .A2(n17108), .B1(
        n17674), .B2(n13840), .ZN(n15779) );
  AOI22_X1 U10158 ( .A1(\pipeline/stageD/target_Jump_temp [7]), .A2(n17676), 
        .B1(n17106), .B2(n15782), .ZN(n15780) );
  AOI22_X1 U10157 ( .A1(\pipeline/data_to_RF_from_WB[7] ), .A2(n17333), .B1(
        \pipeline/Alu_Out_Addr_to_mem[7] ), .B2(n17331), .ZN(n15781) );
  AOI22_X1 U10119 ( .A1(\pipeline/stageF/PC_plus4/N24 ), .A2(n15610), .B1(
        n17674), .B2(n13854), .ZN(n15744) );
  AOI22_X1 U10117 ( .A1(\pipeline/stageD/target_Jump_temp [17]), .A2(n15607), 
        .B1(n17106), .B2(n15747), .ZN(n15745) );
  AOI22_X1 U10116 ( .A1(\pipeline/data_to_RF_from_WB[17] ), .A2(n15605), .B1(
        \pipeline/Alu_Out_Addr_to_mem[17] ), .B2(n15606), .ZN(n15746) );
  AOI22_X1 U10221 ( .A1(\pipeline/stageF/PC_plus4/N8 ), .A2(n17108), .B1(
        n17674), .B2(n13806), .ZN(n15824) );
  AOI22_X1 U10215 ( .A1(\pipeline/stageD/target_Jump_temp [1]), .A2(n17676), 
        .B1(n17106), .B2(n15831), .ZN(n15825) );
  AOI22_X1 U10211 ( .A1(\pipeline/data_to_RF_from_WB[1] ), .A2(n17332), .B1(
        \pipeline/Alu_Out_Addr_to_mem[1] ), .B2(n17330), .ZN(n15826) );
  AOI22_X1 U10184 ( .A1(\pipeline/stageF/PC_plus4/N18 ), .A2(n17108), .B1(
        n17674), .B2(n13824), .ZN(n15799) );
  AOI22_X1 U10182 ( .A1(\pipeline/stageD/target_Jump_temp [11]), .A2(n17675), 
        .B1(n17106), .B2(n15802), .ZN(n15800) );
  AOI22_X1 U10181 ( .A1(\pipeline/data_to_RF_from_WB[11] ), .A2(n17332), .B1(
        \pipeline/Alu_Out_Addr_to_mem[11] ), .B2(n17331), .ZN(n15801) );
  AOI22_X1 U10131 ( .A1(\pipeline/stageF/PC_plus4/N21 ), .A2(n17108), .B1(
        n17674), .B2(n13852), .ZN(n15754) );
  AOI22_X1 U10129 ( .A1(\pipeline/stageD/target_Jump_temp [14]), .A2(n17675), 
        .B1(n17106), .B2(n15757), .ZN(n15755) );
  AOI22_X1 U10128 ( .A1(\pipeline/data_to_RF_from_WB[14] ), .A2(n17333), .B1(
        \pipeline/Alu_Out_Addr_to_mem[14] ), .B2(n17331), .ZN(n15756) );
  AOI22_X1 U10190 ( .A1(\pipeline/stageF/PC_plus4/N16 ), .A2(n17108), .B1(
        n17674), .B2(n13821), .ZN(n15804) );
  AOI22_X1 U10188 ( .A1(\pipeline/stageD/target_Jump_temp [9]), .A2(n15607), 
        .B1(n15608), .B2(n15807), .ZN(n15805) );
  AOI22_X1 U10187 ( .A1(\pipeline/data_to_RF_from_WB[9] ), .A2(n17332), .B1(
        \pipeline/Alu_Out_Addr_to_mem[9] ), .B2(n17331), .ZN(n15806) );
  AOI22_X1 U9967 ( .A1(\pipeline/stageD/offset_jump_sign_ext [24]), .A2(n15600), .B1(n17672), .B2(InstrFetched[24]), .ZN(n15644) );
  AOI22_X1 U9935 ( .A1(n15600), .A2(\pipeline/stageD/offset_to_jump_temp [7]), 
        .B1(n17672), .B2(InstrFetched[7]), .ZN(n15628) );
  AOI22_X1 U9927 ( .A1(n15600), .A2(\pipeline/stageD/offset_to_jump_temp [3]), 
        .B1(n17672), .B2(InstrFetched[3]), .ZN(n15624) );
  AOI22_X1 U9911 ( .A1(n15600), .A2(\pipeline/nextPC_IFID_DEC[16] ), .B1(
        n15601), .B2(\pipeline/stageF/PC_plus4/N23 ), .ZN(n15612) );
  AOI22_X1 U10180 ( .A1(n15600), .A2(\pipeline/nextPC_IFID_DEC[6] ), .B1(
        n15601), .B2(\pipeline/stageF/PC_plus4/N13 ), .ZN(n15798) );
  AOI22_X1 U10085 ( .A1(n15600), .A2(\pipeline/nextPC_IFID_DEC[23] ), .B1(
        n15601), .B2(\pipeline/stageF/PC_plus4/N30 ), .ZN(n15718) );
  AOI21_X1 U9971 ( .B1(InstrFetched[26]), .B2(n15646), .A(n15648), .ZN(n15647)
         );
  OAI21_X1 U9970 ( .B1(n17409), .B2(n15646), .A(n15647), .ZN(n3962) );
  AOI21_X1 U9979 ( .B1(InstrFetched[30]), .B2(n15646), .A(n15648), .ZN(n15652)
         );
  OAI21_X1 U9978 ( .B1(n17347), .B2(n15646), .A(n15652), .ZN(n3958) );
  AOI21_X1 U9975 ( .B1(InstrFetched[28]), .B2(n15646), .A(n15648), .ZN(n15650)
         );
  OAI21_X1 U9974 ( .B1(n17348), .B2(n15646), .A(n15650), .ZN(n3960) );
  NAND2_X1 U10987 ( .A1(n17701), .A2(\pipeline/data_to_RF_from_WB[14] ), .ZN(
        n15094) );
  OAI22_X1 U9555 ( .A1(n17509), .A2(n17418), .B1(n17422), .B2(n15094), .ZN(
        \pipeline/EXMEM_stage/N53 ) );
  NAND2_X1 U10965 ( .A1(n17702), .A2(\pipeline/data_to_RF_from_WB[25] ), .ZN(
        n15072) );
  OAI22_X1 U9532 ( .A1(n17520), .A2(n17418), .B1(n17422), .B2(n15072), .ZN(
        \pipeline/EXMEM_stage/N64 ) );
  NAND2_X1 U10979 ( .A1(n17702), .A2(\pipeline/data_to_RF_from_WB[18] ), .ZN(
        n15086) );
  OAI22_X1 U9547 ( .A1(n17513), .A2(n17418), .B1(n17422), .B2(n15086), .ZN(
        \pipeline/EXMEM_stage/N57 ) );
  NAND2_X1 U10973 ( .A1(n17702), .A2(\pipeline/data_to_RF_from_WB[21] ), .ZN(
        n15080) );
  OAI22_X1 U9540 ( .A1(n17516), .A2(n17418), .B1(n17422), .B2(n15080), .ZN(
        \pipeline/EXMEM_stage/N60 ) );
  NAND2_X1 U10955 ( .A1(n17703), .A2(\pipeline/data_to_RF_from_WB[30] ), .ZN(
        n15062) );
  OAI22_X1 U9522 ( .A1(n17525), .A2(n17418), .B1(n17422), .B2(n15062), .ZN(
        \pipeline/EXMEM_stage/N69 ) );
  NAND2_X1 U10999 ( .A1(n17704), .A2(\pipeline/data_to_RF_from_WB[8] ), .ZN(
        n15106) );
  OAI22_X1 U9569 ( .A1(n17503), .A2(n17418), .B1(n17422), .B2(n15106), .ZN(
        \pipeline/EXMEM_stage/N47 ) );
  NAND2_X1 U10953 ( .A1(n17703), .A2(\pipeline/data_to_RF_from_WB[31] ), .ZN(
        n14988) );
  OAI22_X1 U9487 ( .A1(n17526), .A2(n17418), .B1(n17422), .B2(n14988), .ZN(
        \pipeline/EXMEM_stage/N70 ) );
  NAND2_X1 U11005 ( .A1(n17704), .A2(\pipeline/data_to_RF_from_WB[5] ), .ZN(
        n15112) );
  OAI22_X1 U9575 ( .A1(n17500), .A2(n17418), .B1(n17422), .B2(n15112), .ZN(
        \pipeline/EXMEM_stage/N44 ) );
  NAND2_X1 U11001 ( .A1(n17704), .A2(\pipeline/data_to_RF_from_WB[7] ), .ZN(
        n15108) );
  OAI22_X1 U9571 ( .A1(n17502), .A2(n17418), .B1(n17422), .B2(n15108), .ZN(
        \pipeline/EXMEM_stage/N46 ) );
  NAND2_X1 U11011 ( .A1(n17704), .A2(\pipeline/data_to_RF_from_WB[2] ), .ZN(
        n15118) );
  OAI22_X1 U9581 ( .A1(n17497), .A2(n17418), .B1(n17422), .B2(n15118), .ZN(
        \pipeline/EXMEM_stage/N41 ) );
  NAND2_X1 U10975 ( .A1(n17701), .A2(\pipeline/data_to_RF_from_WB[20] ), .ZN(
        n15082) );
  OAI22_X1 U9543 ( .A1(n17515), .A2(n17418), .B1(n17422), .B2(n15082), .ZN(
        \pipeline/EXMEM_stage/N59 ) );
  NAND2_X1 U10991 ( .A1(n17704), .A2(\pipeline/data_to_RF_from_WB[12] ), .ZN(
        n15098) );
  OAI22_X1 U9559 ( .A1(n17507), .A2(n17418), .B1(n17422), .B2(n15098), .ZN(
        \pipeline/EXMEM_stage/N51 ) );
  NAND2_X1 U10985 ( .A1(n17702), .A2(\pipeline/data_to_RF_from_WB[15] ), .ZN(
        n15092) );
  OAI22_X1 U9553 ( .A1(n17510), .A2(n17418), .B1(n17422), .B2(n15092), .ZN(
        \pipeline/EXMEM_stage/N54 ) );
  NAND2_X1 U10995 ( .A1(n17704), .A2(\pipeline/data_to_RF_from_WB[10] ), .ZN(
        n15102) );
  OAI22_X1 U9565 ( .A1(n17505), .A2(n17418), .B1(n17422), .B2(n15102), .ZN(
        \pipeline/EXMEM_stage/N49 ) );
  NAND2_X1 U10997 ( .A1(n17704), .A2(\pipeline/data_to_RF_from_WB[9] ), .ZN(
        n15104) );
  OAI22_X1 U9567 ( .A1(n17504), .A2(n17418), .B1(n17422), .B2(n15104), .ZN(
        \pipeline/EXMEM_stage/N48 ) );
  NAND2_X1 U10981 ( .A1(n17701), .A2(\pipeline/data_to_RF_from_WB[17] ), .ZN(
        n15088) );
  OAI22_X1 U9549 ( .A1(n17512), .A2(n17418), .B1(n17422), .B2(n15088), .ZN(
        \pipeline/EXMEM_stage/N56 ) );
  NAND2_X1 U10969 ( .A1(n17701), .A2(\pipeline/data_to_RF_from_WB[23] ), .ZN(
        n15076) );
  OAI22_X1 U9536 ( .A1(n17518), .A2(n17418), .B1(n17422), .B2(n15076), .ZN(
        \pipeline/EXMEM_stage/N62 ) );
  NAND2_X1 U10983 ( .A1(n17702), .A2(\pipeline/data_to_RF_from_WB[16] ), .ZN(
        n15090) );
  OAI22_X1 U9551 ( .A1(n17511), .A2(n17418), .B1(n17422), .B2(n15090), .ZN(
        \pipeline/EXMEM_stage/N55 ) );
  NAND2_X1 U10977 ( .A1(n17701), .A2(\pipeline/data_to_RF_from_WB[19] ), .ZN(
        n15084) );
  OAI22_X1 U9545 ( .A1(n17514), .A2(n17418), .B1(n17422), .B2(n15084), .ZN(
        \pipeline/EXMEM_stage/N58 ) );
  NAND2_X1 U10963 ( .A1(n17702), .A2(\pipeline/data_to_RF_from_WB[26] ), .ZN(
        n15070) );
  OAI22_X1 U9530 ( .A1(n17521), .A2(n17418), .B1(n17422), .B2(n15070), .ZN(
        \pipeline/EXMEM_stage/N65 ) );
  NAND2_X1 U11007 ( .A1(n17704), .A2(\pipeline/data_to_RF_from_WB[4] ), .ZN(
        n15114) );
  OAI22_X1 U9577 ( .A1(n17499), .A2(n17418), .B1(n17422), .B2(n15114), .ZN(
        \pipeline/EXMEM_stage/N43 ) );
  NAND2_X1 U10989 ( .A1(n17704), .A2(\pipeline/data_to_RF_from_WB[13] ), .ZN(
        n15096) );
  OAI22_X1 U9557 ( .A1(n17508), .A2(n17418), .B1(n17422), .B2(n15096), .ZN(
        \pipeline/EXMEM_stage/N52 ) );
  NAND2_X1 U10959 ( .A1(n17703), .A2(\pipeline/data_to_RF_from_WB[28] ), .ZN(
        n15066) );
  OAI22_X1 U9526 ( .A1(n17523), .A2(n17418), .B1(n17422), .B2(n15066), .ZN(
        \pipeline/EXMEM_stage/N67 ) );
  NAND2_X1 U10967 ( .A1(n17701), .A2(\pipeline/data_to_RF_from_WB[24] ), .ZN(
        n15074) );
  OAI22_X1 U9534 ( .A1(n17519), .A2(n17418), .B1(n17422), .B2(n15074), .ZN(
        \pipeline/EXMEM_stage/N63 ) );
  NAND2_X1 U10971 ( .A1(n17701), .A2(\pipeline/data_to_RF_from_WB[22] ), .ZN(
        n15078) );
  OAI22_X1 U9538 ( .A1(n17517), .A2(n17418), .B1(n17422), .B2(n15078), .ZN(
        \pipeline/EXMEM_stage/N61 ) );
  NAND2_X1 U11003 ( .A1(n17704), .A2(\pipeline/data_to_RF_from_WB[6] ), .ZN(
        n15110) );
  OAI22_X1 U9573 ( .A1(n17501), .A2(n17418), .B1(n17422), .B2(n15110), .ZN(
        \pipeline/EXMEM_stage/N45 ) );
  NAND2_X1 U11013 ( .A1(n17704), .A2(\pipeline/data_to_RF_from_WB[1] ), .ZN(
        n15120) );
  OAI22_X1 U9583 ( .A1(n17496), .A2(n17418), .B1(n17422), .B2(n15120), .ZN(
        \pipeline/EXMEM_stage/N40 ) );
  NAND2_X1 U10957 ( .A1(n17703), .A2(\pipeline/data_to_RF_from_WB[29] ), .ZN(
        n15064) );
  OAI22_X1 U9524 ( .A1(n17524), .A2(n17418), .B1(n17422), .B2(n15064), .ZN(
        \pipeline/EXMEM_stage/N68 ) );
  NAND2_X1 U11015 ( .A1(n17704), .A2(\pipeline/data_to_RF_from_WB[0] ), .ZN(
        n15122) );
  OAI22_X1 U9587 ( .A1(n17495), .A2(n17418), .B1(n17422), .B2(n15122), .ZN(
        \pipeline/EXMEM_stage/N39 ) );
  NAND2_X1 U10961 ( .A1(n17703), .A2(\pipeline/data_to_RF_from_WB[27] ), .ZN(
        n15068) );
  OAI22_X1 U9528 ( .A1(n17522), .A2(n17418), .B1(n17422), .B2(n15068), .ZN(
        \pipeline/EXMEM_stage/N66 ) );
  NAND2_X1 U11009 ( .A1(n17703), .A2(\pipeline/data_to_RF_from_WB[3] ), .ZN(
        n15116) );
  OAI22_X1 U9579 ( .A1(n17498), .A2(n17418), .B1(n17422), .B2(n15116), .ZN(
        \pipeline/EXMEM_stage/N42 ) );
  NAND2_X1 U10993 ( .A1(n17704), .A2(\pipeline/data_to_RF_from_WB[11] ), .ZN(
        n15100) );
  OAI22_X1 U9561 ( .A1(n17506), .A2(n17418), .B1(n17422), .B2(n15100), .ZN(
        \pipeline/EXMEM_stage/N50 ) );
  NOR2_X1 U8678 ( .A1(n17431), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N181 ) );
  AOI22_X1 U8989 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[31][18] ), .A2(n17154), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[30][18] ), .B2(n17683), .ZN(
        n14508) );
  AOI22_X1 U8988 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[29][18] ), .A2(n17684), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[28][18] ), .B2(n17685), .ZN(
        n14509) );
  NAND2_X1 U9375 ( .A1(n17408), .A2(n17329), .ZN(n14860) );
  AOI222_X1 U8987 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[4][18] ), .A2(n17686), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[25][18] ), .B2(n17153), .C1(
        \pipeline/RegFile_DEC_WB/RegBank[24][18] ), .C2(n17687), .ZN(n14510)
         );
  AOI22_X1 U8986 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[27][18] ), .A2(n17688), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[26][18] ), .B2(n17689), .ZN(
        n14504) );
  AOI22_X1 U8985 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[23][18] ), .A2(n17690), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[22][18] ), .B2(n17691), .ZN(
        n14505) );
  AOI22_X1 U8984 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[21][18] ), .A2(n17692), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[20][18] ), .B2(n17693), .ZN(
        n14506) );
  AOI22_X1 U8983 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[19][18] ), .A2(n17694), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[18][18] ), .B2(n17695), .ZN(
        n14507) );
  NAND4_X1 U8982 ( .A1(n14504), .A2(n14505), .A3(n14506), .A4(n14507), .ZN(
        n14493) );
  AOI22_X1 U8981 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[17][18] ), .A2(n17696), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[16][18] ), .B2(n17697), .ZN(
        n14500) );
  NOR2_X1 U9353 ( .A1(n14865), .A2(n14867), .ZN(n14226) );
  AOI22_X1 U8980 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[12][18] ), .A2(n17698), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[13][18] ), .B2(n14226), .ZN(
        n14501) );
  AOI22_X1 U8979 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[8][18] ), .A2(n14223), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[15][18] ), .B2(n17152), .ZN(
        n14502) );
  NOR2_X1 U9348 ( .A1(n14860), .A2(n14867), .ZN(n14221) );
  AOI22_X1 U8978 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[9][18] ), .A2(n14221), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[10][18] ), .B2(n17699), .ZN(
        n14503) );
  NAND4_X1 U8977 ( .A1(n14500), .A2(n14501), .A3(n14502), .A4(n14503), .ZN(
        n14494) );
  AOI22_X1 U8976 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[11][18] ), .A2(n17151), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[3][18] ), .B2(n14216), .ZN(n14496) );
  AOI22_X1 U8975 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[14][18] ), .A2(n17700), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[5][18] ), .B2(n14214), .ZN(n14497) );
  AOI22_X1 U8974 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[2][18] ), .A2(n17367), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[7][18] ), .B2(n14212), .ZN(n14498) );
  AOI22_X1 U8973 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[6][18] ), .A2(n17368), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[1][18] ), .B2(n14210), .ZN(n14499) );
  NAND4_X1 U8972 ( .A1(n14496), .A2(n14497), .A3(n14498), .A4(n14499), .ZN(
        n14495) );
  NOR4_X1 U8971 ( .A1(n14492), .A2(n14493), .A3(n14494), .A4(n14495), .ZN(
        n14491) );
  NOR2_X1 U8970 ( .A1(n14491), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N152 ) );
  AOI22_X1 U9229 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[31][6] ), .A2(n17154), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[30][6] ), .B2(n17683), .ZN(n14748) );
  AOI22_X1 U9228 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[29][6] ), .A2(n17684), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[28][6] ), .B2(n17685), .ZN(n14749) );
  AOI222_X1 U9227 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[4][6] ), .A2(n17686), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[25][6] ), .B2(n17153), .C1(
        \pipeline/RegFile_DEC_WB/RegBank[24][6] ), .C2(n17687), .ZN(n14750) );
  AOI22_X1 U9226 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[27][6] ), .A2(n17688), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[26][6] ), .B2(n17689), .ZN(n14744) );
  AOI22_X1 U9225 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[23][6] ), .A2(n17690), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[22][6] ), .B2(n17691), .ZN(n14745) );
  AOI22_X1 U9224 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[21][6] ), .A2(n17692), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[20][6] ), .B2(n17693), .ZN(n14746) );
  AOI22_X1 U9223 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[19][6] ), .A2(n17694), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[18][6] ), .B2(n17695), .ZN(n14747) );
  NAND4_X1 U9222 ( .A1(n14744), .A2(n14745), .A3(n14746), .A4(n14747), .ZN(
        n14733) );
  AOI22_X1 U9221 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[17][6] ), .A2(n17696), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[16][6] ), .B2(n17697), .ZN(n14740) );
  AOI22_X1 U9220 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[12][6] ), .A2(n17698), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[13][6] ), .B2(n17358), .ZN(n14741) );
  AOI22_X1 U9219 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[8][6] ), .A2(n17417), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[15][6] ), .B2(n17152), .ZN(n14742) );
  AOI22_X1 U9218 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[9][6] ), .A2(n17352), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[10][6] ), .B2(n17699), .ZN(n14743) );
  NAND4_X1 U9217 ( .A1(n14740), .A2(n14741), .A3(n14742), .A4(n14743), .ZN(
        n14734) );
  AOI22_X1 U9216 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[11][6] ), .A2(n17151), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[3][6] ), .B2(n17413), .ZN(n14736)
         );
  AOI22_X1 U9215 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[14][6] ), .A2(n17700), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[5][6] ), .B2(n17414), .ZN(n14737)
         );
  AOI22_X1 U9214 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[2][6] ), .A2(n17355), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[7][6] ), .B2(n17415), .ZN(n14738)
         );
  AOI22_X1 U9213 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[6][6] ), .A2(n17356), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[1][6] ), .B2(n17416), .ZN(n14739)
         );
  NAND4_X1 U9212 ( .A1(n14736), .A2(n14737), .A3(n14738), .A4(n14739), .ZN(
        n14735) );
  NOR4_X1 U9211 ( .A1(n14732), .A2(n14733), .A3(n14734), .A4(n14735), .ZN(
        n14731) );
  NOR2_X1 U9210 ( .A1(n14731), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N140 ) );
  AOI22_X1 U9169 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[31][9] ), .A2(n17154), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[30][9] ), .B2(n17683), .ZN(n14688) );
  AOI22_X1 U9168 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[29][9] ), .A2(n17684), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[28][9] ), .B2(n17685), .ZN(n14689) );
  AOI222_X1 U9167 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[4][9] ), .A2(n17686), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[25][9] ), .B2(n17153), .C1(
        \pipeline/RegFile_DEC_WB/RegBank[24][9] ), .C2(n14246), .ZN(n14690) );
  AOI22_X1 U9166 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[27][9] ), .A2(n17688), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[26][9] ), .B2(n17689), .ZN(n14684) );
  AOI22_X1 U9165 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[23][9] ), .A2(n17690), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[22][9] ), .B2(n17691), .ZN(n14685) );
  AOI22_X1 U9164 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[21][9] ), .A2(n17692), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[20][9] ), .B2(n17693), .ZN(n14686) );
  AOI22_X1 U9163 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[19][9] ), .A2(n17694), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[18][9] ), .B2(n17695), .ZN(n14687) );
  NAND4_X1 U9162 ( .A1(n14684), .A2(n14685), .A3(n14686), .A4(n14687), .ZN(
        n14673) );
  AOI22_X1 U9161 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[17][9] ), .A2(n17696), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[16][9] ), .B2(n17697), .ZN(n14680) );
  AOI22_X1 U9160 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[12][9] ), .A2(n17698), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[13][9] ), .B2(n17358), .ZN(n14681) );
  AOI22_X1 U9159 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[8][9] ), .A2(n14223), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[15][9] ), .B2(n17152), .ZN(n14682) );
  AOI22_X1 U9158 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[9][9] ), .A2(n17352), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[10][9] ), .B2(n17699), .ZN(n14683) );
  NAND4_X1 U9157 ( .A1(n14680), .A2(n14681), .A3(n14682), .A4(n14683), .ZN(
        n14674) );
  AOI22_X1 U9156 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[11][9] ), .A2(n17151), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[3][9] ), .B2(n14216), .ZN(n14676)
         );
  AOI22_X1 U9155 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[14][9] ), .A2(n17700), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[5][9] ), .B2(n14214), .ZN(n14677)
         );
  AOI22_X1 U9154 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[2][9] ), .A2(n17355), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[7][9] ), .B2(n14212), .ZN(n14678)
         );
  AOI22_X1 U9153 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[6][9] ), .A2(n17356), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[1][9] ), .B2(n14210), .ZN(n14679)
         );
  NAND4_X1 U9152 ( .A1(n14676), .A2(n14677), .A3(n14678), .A4(n14679), .ZN(
        n14675) );
  NOR4_X1 U9151 ( .A1(n14672), .A2(n14673), .A3(n14674), .A4(n14675), .ZN(
        n14671) );
  NOR2_X1 U9150 ( .A1(n14671), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N143 ) );
  AOI22_X1 U8809 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[31][27] ), .A2(n14249), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[30][27] ), .B2(n14250), .ZN(
        n14328) );
  AOI22_X1 U8808 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[29][27] ), .A2(n14247), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[28][27] ), .B2(n14248), .ZN(
        n14329) );
  AOI222_X1 U8807 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[4][27] ), .A2(n14244), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[25][27] ), .B2(n14245), .C1(
        \pipeline/RegFile_DEC_WB/RegBank[24][27] ), .C2(n17687), .ZN(n14330)
         );
  AOI22_X1 U8806 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[27][27] ), .A2(n14239), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[26][27] ), .B2(n14240), .ZN(
        n14324) );
  AOI22_X1 U8805 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[23][27] ), .A2(n14237), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[22][27] ), .B2(n14238), .ZN(
        n14325) );
  AOI22_X1 U8804 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[21][27] ), .A2(n14235), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[20][27] ), .B2(n14236), .ZN(
        n14326) );
  AOI22_X1 U8803 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[19][27] ), .A2(n14233), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[18][27] ), .B2(n14234), .ZN(
        n14327) );
  NAND4_X1 U8802 ( .A1(n14324), .A2(n14325), .A3(n14326), .A4(n14327), .ZN(
        n14313) );
  AOI22_X1 U8801 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[17][27] ), .A2(n14227), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[16][27] ), .B2(n14228), .ZN(
        n14320) );
  AOI22_X1 U8800 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[12][27] ), .A2(n14225), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[13][27] ), .B2(n17357), .ZN(
        n14321) );
  AOI22_X1 U8799 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[8][27] ), .A2(n17417), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[15][27] ), .B2(n17152), .ZN(
        n14322) );
  AOI22_X1 U8798 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[9][27] ), .A2(n17351), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[10][27] ), .B2(n14222), .ZN(
        n14323) );
  NAND4_X1 U8797 ( .A1(n14320), .A2(n14321), .A3(n14322), .A4(n14323), .ZN(
        n14314) );
  AOI22_X1 U8796 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[11][27] ), .A2(n17151), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[3][27] ), .B2(n17413), .ZN(n14316) );
  AOI22_X1 U8795 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[14][27] ), .A2(n17700), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[5][27] ), .B2(n17414), .ZN(n14317) );
  AOI22_X1 U8794 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[2][27] ), .A2(n17353), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[7][27] ), .B2(n17415), .ZN(n14318) );
  AOI22_X1 U8793 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[6][27] ), .A2(n17354), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[1][27] ), .B2(n17416), .ZN(n14319) );
  NAND4_X1 U8792 ( .A1(n14316), .A2(n14317), .A3(n14318), .A4(n14319), .ZN(
        n14315) );
  NOR4_X1 U8791 ( .A1(n14312), .A2(n14313), .A3(n14314), .A4(n14315), .ZN(
        n14311) );
  NOR2_X1 U8790 ( .A1(n14311), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N161 ) );
  AOI22_X1 U8969 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[31][19] ), .A2(n17154), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[30][19] ), .B2(n17683), .ZN(
        n14488) );
  AOI22_X1 U8968 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[29][19] ), .A2(n17684), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[28][19] ), .B2(n17685), .ZN(
        n14489) );
  AOI222_X1 U8967 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[4][19] ), .A2(n17686), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[25][19] ), .B2(n17153), .C1(
        \pipeline/RegFile_DEC_WB/RegBank[24][19] ), .C2(n17687), .ZN(n14490)
         );
  AOI22_X1 U8966 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[27][19] ), .A2(n17688), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[26][19] ), .B2(n17689), .ZN(
        n14484) );
  AOI22_X1 U8965 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[23][19] ), .A2(n17690), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[22][19] ), .B2(n17691), .ZN(
        n14485) );
  AOI22_X1 U8964 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[21][19] ), .A2(n17692), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[20][19] ), .B2(n17693), .ZN(
        n14486) );
  AOI22_X1 U8963 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[19][19] ), .A2(n17694), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[18][19] ), .B2(n17695), .ZN(
        n14487) );
  NAND4_X1 U8962 ( .A1(n14484), .A2(n14485), .A3(n14486), .A4(n14487), .ZN(
        n14473) );
  AOI22_X1 U8961 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[17][19] ), .A2(n17696), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[16][19] ), .B2(n17697), .ZN(
        n14480) );
  AOI22_X1 U8960 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[12][19] ), .A2(n17698), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[13][19] ), .B2(n14226), .ZN(
        n14481) );
  AOI22_X1 U8959 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[8][19] ), .A2(n14223), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[15][19] ), .B2(n17152), .ZN(
        n14482) );
  AOI22_X1 U8958 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[9][19] ), .A2(n14221), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[10][19] ), .B2(n17699), .ZN(
        n14483) );
  NAND4_X1 U8957 ( .A1(n14480), .A2(n14481), .A3(n14482), .A4(n14483), .ZN(
        n14474) );
  AOI22_X1 U8956 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[11][19] ), .A2(n17151), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[3][19] ), .B2(n14216), .ZN(n14476) );
  AOI22_X1 U8955 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[14][19] ), .A2(n17700), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[5][19] ), .B2(n14214), .ZN(n14477) );
  AOI22_X1 U8954 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[2][19] ), .A2(n17367), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[7][19] ), .B2(n14212), .ZN(n14478) );
  AOI22_X1 U8953 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[6][19] ), .A2(n17368), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[1][19] ), .B2(n14210), .ZN(n14479) );
  NAND4_X1 U8952 ( .A1(n14476), .A2(n14477), .A3(n14478), .A4(n14479), .ZN(
        n14475) );
  NOR4_X1 U8951 ( .A1(n14472), .A2(n14473), .A3(n14474), .A4(n14475), .ZN(
        n14471) );
  NOR2_X1 U8950 ( .A1(n14471), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N153 ) );
  AOI22_X1 U9049 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[31][15] ), .A2(n17154), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[30][15] ), .B2(n17683), .ZN(
        n14568) );
  AOI22_X1 U9048 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[29][15] ), .A2(n17684), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[28][15] ), .B2(n17685), .ZN(
        n14569) );
  AOI222_X1 U9047 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[4][15] ), .A2(n17686), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[25][15] ), .B2(n17153), .C1(
        \pipeline/RegFile_DEC_WB/RegBank[24][15] ), .C2(n17687), .ZN(n14570)
         );
  AOI22_X1 U9046 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[27][15] ), .A2(n17688), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[26][15] ), .B2(n17689), .ZN(
        n14564) );
  AOI22_X1 U9045 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[23][15] ), .A2(n17690), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[22][15] ), .B2(n17691), .ZN(
        n14565) );
  AOI22_X1 U9044 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[21][15] ), .A2(n17692), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[20][15] ), .B2(n17693), .ZN(
        n14566) );
  AOI22_X1 U9043 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[19][15] ), .A2(n17694), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[18][15] ), .B2(n17695), .ZN(
        n14567) );
  NAND4_X1 U9042 ( .A1(n14564), .A2(n14565), .A3(n14566), .A4(n14567), .ZN(
        n14553) );
  AOI22_X1 U9041 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[17][15] ), .A2(n17696), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[16][15] ), .B2(n17697), .ZN(
        n14560) );
  AOI22_X1 U9040 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[12][15] ), .A2(n17698), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[13][15] ), .B2(n17358), .ZN(
        n14561) );
  AOI22_X1 U9039 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[8][15] ), .A2(n14223), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[15][15] ), .B2(n17152), .ZN(
        n14562) );
  AOI22_X1 U9038 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[9][15] ), .A2(n17352), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[10][15] ), .B2(n17699), .ZN(
        n14563) );
  NAND4_X1 U9037 ( .A1(n14560), .A2(n14561), .A3(n14562), .A4(n14563), .ZN(
        n14554) );
  AOI22_X1 U9036 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[11][15] ), .A2(n17151), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[3][15] ), .B2(n14216), .ZN(n14556) );
  AOI22_X1 U9035 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[14][15] ), .A2(n17700), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[5][15] ), .B2(n14214), .ZN(n14557) );
  AOI22_X1 U9034 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[2][15] ), .A2(n17355), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[7][15] ), .B2(n14212), .ZN(n14558) );
  AOI22_X1 U9033 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[6][15] ), .A2(n17356), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[1][15] ), .B2(n14210), .ZN(n14559) );
  NAND4_X1 U9032 ( .A1(n14556), .A2(n14557), .A3(n14558), .A4(n14559), .ZN(
        n14555) );
  NOR4_X1 U9031 ( .A1(n14552), .A2(n14553), .A3(n14554), .A4(n14555), .ZN(
        n14551) );
  NOR2_X1 U9030 ( .A1(n14551), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N149 ) );
  AOI22_X1 U9009 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[31][17] ), .A2(n17154), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[30][17] ), .B2(n17683), .ZN(
        n14528) );
  AOI22_X1 U9008 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[29][17] ), .A2(n17684), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[28][17] ), .B2(n17685), .ZN(
        n14529) );
  AOI222_X1 U9007 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[4][17] ), .A2(n17686), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[25][17] ), .B2(n17153), .C1(
        \pipeline/RegFile_DEC_WB/RegBank[24][17] ), .C2(n17687), .ZN(n14530)
         );
  AOI22_X1 U9006 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[27][17] ), .A2(n17688), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[26][17] ), .B2(n17689), .ZN(
        n14524) );
  AOI22_X1 U9005 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[23][17] ), .A2(n17690), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[22][17] ), .B2(n17691), .ZN(
        n14525) );
  AOI22_X1 U9004 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[21][17] ), .A2(n17692), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[20][17] ), .B2(n17693), .ZN(
        n14526) );
  AOI22_X1 U9003 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[19][17] ), .A2(n17694), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[18][17] ), .B2(n17695), .ZN(
        n14527) );
  NAND4_X1 U9002 ( .A1(n14524), .A2(n14525), .A3(n14526), .A4(n14527), .ZN(
        n14513) );
  AOI22_X1 U9001 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[17][17] ), .A2(n17696), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[16][17] ), .B2(n17697), .ZN(
        n14520) );
  AOI22_X1 U9000 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[12][17] ), .A2(n17698), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[13][17] ), .B2(n14226), .ZN(
        n14521) );
  AOI22_X1 U8999 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[8][17] ), .A2(n14223), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[15][17] ), .B2(n17152), .ZN(
        n14522) );
  AOI22_X1 U8998 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[9][17] ), .A2(n14221), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[10][17] ), .B2(n17699), .ZN(
        n14523) );
  NAND4_X1 U8997 ( .A1(n14520), .A2(n14521), .A3(n14522), .A4(n14523), .ZN(
        n14514) );
  AOI22_X1 U8996 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[11][17] ), .A2(n17151), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[3][17] ), .B2(n14216), .ZN(n14516) );
  AOI22_X1 U8995 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[14][17] ), .A2(n17700), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[5][17] ), .B2(n14214), .ZN(n14517) );
  AOI22_X1 U8994 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[2][17] ), .A2(n17367), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[7][17] ), .B2(n14212), .ZN(n14518) );
  AOI22_X1 U8993 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[6][17] ), .A2(n17368), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[1][17] ), .B2(n14210), .ZN(n14519) );
  NAND4_X1 U8992 ( .A1(n14516), .A2(n14517), .A3(n14518), .A4(n14519), .ZN(
        n14515) );
  NOR4_X1 U8991 ( .A1(n14512), .A2(n14513), .A3(n14514), .A4(n14515), .ZN(
        n14511) );
  NOR2_X1 U8990 ( .A1(n14511), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N151 ) );
  AOI22_X1 U9385 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[31][0] ), .A2(n14249), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[30][0] ), .B2(n14250), .ZN(n14880) );
  AOI22_X1 U9380 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[29][0] ), .A2(n14247), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[28][0] ), .B2(n14248), .ZN(n14881) );
  AOI222_X1 U9372 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[4][0] ), .A2(n14244), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[25][0] ), .B2(n17153), .C1(
        \pipeline/RegFile_DEC_WB/RegBank[24][0] ), .C2(n17687), .ZN(n14882) );
  AOI22_X1 U9368 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[27][0] ), .A2(n14239), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[26][0] ), .B2(n14240), .ZN(n14874) );
  AOI22_X1 U9365 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[23][0] ), .A2(n14237), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[22][0] ), .B2(n14238), .ZN(n14875) );
  AOI22_X1 U9362 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[21][0] ), .A2(n14235), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[20][0] ), .B2(n14236), .ZN(n14876) );
  AOI22_X1 U9359 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[19][0] ), .A2(n14233), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[18][0] ), .B2(n14234), .ZN(n14877) );
  NAND4_X1 U9358 ( .A1(n14874), .A2(n14875), .A3(n14876), .A4(n14877), .ZN(
        n14853) );
  AOI22_X1 U9355 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[17][0] ), .A2(n14227), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[16][0] ), .B2(n14228), .ZN(n14868) );
  AOI22_X1 U9352 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[12][0] ), .A2(n14225), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[13][0] ), .B2(n17357), .ZN(n14869) );
  AOI22_X1 U9349 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[8][0] ), .A2(n17417), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[15][0] ), .B2(n17152), .ZN(n14870) );
  AOI22_X1 U9346 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[9][0] ), .A2(n17351), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[10][0] ), .B2(n14222), .ZN(n14871) );
  NAND4_X1 U9345 ( .A1(n14868), .A2(n14869), .A3(n14870), .A4(n14871), .ZN(
        n14854) );
  AOI22_X1 U9342 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[11][0] ), .A2(n17151), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[3][0] ), .B2(n17413), .ZN(n14856)
         );
  AOI22_X1 U9339 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[14][0] ), .A2(n17700), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[5][0] ), .B2(n17414), .ZN(n14857)
         );
  AOI22_X1 U9336 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[2][0] ), .A2(n17353), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[7][0] ), .B2(n17415), .ZN(n14858)
         );
  AOI22_X1 U9333 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[6][0] ), .A2(n17354), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[1][0] ), .B2(n17416), .ZN(n14859)
         );
  NAND4_X1 U9332 ( .A1(n14856), .A2(n14857), .A3(n14858), .A4(n14859), .ZN(
        n14855) );
  NOR4_X1 U9331 ( .A1(n14852), .A2(n14853), .A3(n14854), .A4(n14855), .ZN(
        n14851) );
  NOR2_X1 U9330 ( .A1(n14851), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N134 ) );
  AOI22_X1 U9269 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[31][4] ), .A2(n17154), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[30][4] ), .B2(n17683), .ZN(n14788) );
  AOI22_X1 U9268 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[29][4] ), .A2(n17684), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[28][4] ), .B2(n17685), .ZN(n14789) );
  AOI222_X1 U9267 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[4][4] ), .A2(n17686), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[25][4] ), .B2(n17153), .C1(
        \pipeline/RegFile_DEC_WB/RegBank[24][4] ), .C2(n14246), .ZN(n14790) );
  AOI22_X1 U9266 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[27][4] ), .A2(n17688), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[26][4] ), .B2(n17689), .ZN(n14784) );
  AOI22_X1 U9265 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[23][4] ), .A2(n17690), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[22][4] ), .B2(n17691), .ZN(n14785) );
  AOI22_X1 U9264 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[21][4] ), .A2(n17692), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[20][4] ), .B2(n17693), .ZN(n14786) );
  AOI22_X1 U9263 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[19][4] ), .A2(n17694), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[18][4] ), .B2(n17695), .ZN(n14787) );
  NAND4_X1 U9262 ( .A1(n14784), .A2(n14785), .A3(n14786), .A4(n14787), .ZN(
        n14773) );
  AOI22_X1 U9261 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[17][4] ), .A2(n17696), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[16][4] ), .B2(n17697), .ZN(n14780) );
  AOI22_X1 U9260 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[12][4] ), .A2(n17698), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[13][4] ), .B2(n17357), .ZN(n14781) );
  AOI22_X1 U9259 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[8][4] ), .A2(n17417), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[15][4] ), .B2(n17152), .ZN(n14782) );
  AOI22_X1 U9258 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[9][4] ), .A2(n17351), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[10][4] ), .B2(n17699), .ZN(n14783) );
  NAND4_X1 U9257 ( .A1(n14780), .A2(n14781), .A3(n14782), .A4(n14783), .ZN(
        n14774) );
  AOI22_X1 U9256 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[11][4] ), .A2(n14215), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[3][4] ), .B2(n17413), .ZN(n14776)
         );
  AOI22_X1 U9255 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[14][4] ), .A2(n17700), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[5][4] ), .B2(n17414), .ZN(n14777)
         );
  AOI22_X1 U9254 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[2][4] ), .A2(n17353), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[7][4] ), .B2(n17415), .ZN(n14778)
         );
  AOI22_X1 U9253 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[6][4] ), .A2(n17354), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[1][4] ), .B2(n17416), .ZN(n14779)
         );
  NAND4_X1 U9252 ( .A1(n14776), .A2(n14777), .A3(n14778), .A4(n14779), .ZN(
        n14775) );
  NOR4_X1 U9251 ( .A1(n14772), .A2(n14773), .A3(n14774), .A4(n14775), .ZN(
        n14771) );
  NOR2_X1 U9250 ( .A1(n14771), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N138 ) );
  AOI22_X1 U8909 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[31][22] ), .A2(n17154), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[30][22] ), .B2(n17683), .ZN(
        n14428) );
  AOI22_X1 U8908 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[29][22] ), .A2(n17684), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[28][22] ), .B2(n17685), .ZN(
        n14429) );
  AOI222_X1 U8907 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[4][22] ), .A2(n17686), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[25][22] ), .B2(n14245), .C1(
        \pipeline/RegFile_DEC_WB/RegBank[24][22] ), .C2(n14246), .ZN(n14430)
         );
  AOI22_X1 U8906 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[27][22] ), .A2(n14239), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[26][22] ), .B2(n17689), .ZN(
        n14424) );
  AOI22_X1 U8905 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[23][22] ), .A2(n17690), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[22][22] ), .B2(n17691), .ZN(
        n14425) );
  AOI22_X1 U8904 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[21][22] ), .A2(n14235), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[20][22] ), .B2(n17693), .ZN(
        n14426) );
  AOI22_X1 U8903 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[19][22] ), .A2(n17694), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[18][22] ), .B2(n17695), .ZN(
        n14427) );
  NAND4_X1 U8902 ( .A1(n14424), .A2(n14425), .A3(n14426), .A4(n14427), .ZN(
        n14413) );
  AOI22_X1 U8901 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[17][22] ), .A2(n14227), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[16][22] ), .B2(n17697), .ZN(
        n14420) );
  AOI22_X1 U8900 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[12][22] ), .A2(n17698), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[13][22] ), .B2(n17357), .ZN(
        n14421) );
  AOI22_X1 U8899 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[8][22] ), .A2(n17417), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[15][22] ), .B2(n17152), .ZN(
        n14422) );
  AOI22_X1 U8898 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[9][22] ), .A2(n17351), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[10][22] ), .B2(n17699), .ZN(
        n14423) );
  NAND4_X1 U8897 ( .A1(n14420), .A2(n14421), .A3(n14422), .A4(n14423), .ZN(
        n14414) );
  AOI22_X1 U8896 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[11][22] ), .A2(n14215), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[3][22] ), .B2(n17413), .ZN(n14416) );
  AOI22_X1 U8895 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[14][22] ), .A2(n14213), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[5][22] ), .B2(n17414), .ZN(n14417) );
  AOI22_X1 U8894 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[2][22] ), .A2(n17353), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[7][22] ), .B2(n17415), .ZN(n14418) );
  AOI22_X1 U8893 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[6][22] ), .A2(n17354), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[1][22] ), .B2(n17416), .ZN(n14419) );
  NAND4_X1 U8892 ( .A1(n14416), .A2(n14417), .A3(n14418), .A4(n14419), .ZN(
        n14415) );
  NOR4_X1 U8891 ( .A1(n14412), .A2(n14413), .A3(n14414), .A4(n14415), .ZN(
        n14411) );
  NOR2_X1 U8890 ( .A1(n14411), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N156 ) );
  AOI22_X1 U9249 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[31][5] ), .A2(n17154), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[30][5] ), .B2(n17683), .ZN(n14768) );
  AOI22_X1 U9248 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[29][5] ), .A2(n17684), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[28][5] ), .B2(n17685), .ZN(n14769) );
  AOI222_X1 U9247 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[4][5] ), .A2(n17686), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[25][5] ), .B2(n17153), .C1(
        \pipeline/RegFile_DEC_WB/RegBank[24][5] ), .C2(n17687), .ZN(n14770) );
  AOI22_X1 U9246 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[27][5] ), .A2(n17688), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[26][5] ), .B2(n17689), .ZN(n14764) );
  AOI22_X1 U9245 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[23][5] ), .A2(n17690), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[22][5] ), .B2(n17691), .ZN(n14765) );
  AOI22_X1 U9244 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[21][5] ), .A2(n17692), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[20][5] ), .B2(n17693), .ZN(n14766) );
  AOI22_X1 U9243 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[19][5] ), .A2(n17694), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[18][5] ), .B2(n17695), .ZN(n14767) );
  NAND4_X1 U9242 ( .A1(n14764), .A2(n14765), .A3(n14766), .A4(n14767), .ZN(
        n14753) );
  AOI22_X1 U9241 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[17][5] ), .A2(n17696), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[16][5] ), .B2(n17697), .ZN(n14760) );
  AOI22_X1 U9240 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[12][5] ), .A2(n17698), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[13][5] ), .B2(n17357), .ZN(n14761) );
  AOI22_X1 U9239 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[8][5] ), .A2(n17417), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[15][5] ), .B2(n17152), .ZN(n14762) );
  AOI22_X1 U9238 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[9][5] ), .A2(n17351), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[10][5] ), .B2(n17699), .ZN(n14763) );
  NAND4_X1 U9237 ( .A1(n14760), .A2(n14761), .A3(n14762), .A4(n14763), .ZN(
        n14754) );
  AOI22_X1 U9236 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[11][5] ), .A2(n14215), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[3][5] ), .B2(n17413), .ZN(n14756)
         );
  AOI22_X1 U9235 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[14][5] ), .A2(n17700), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[5][5] ), .B2(n17414), .ZN(n14757)
         );
  AOI22_X1 U9234 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[2][5] ), .A2(n17353), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[7][5] ), .B2(n17415), .ZN(n14758)
         );
  AOI22_X1 U9233 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[6][5] ), .A2(n17354), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[1][5] ), .B2(n17416), .ZN(n14759)
         );
  NAND4_X1 U9232 ( .A1(n14756), .A2(n14757), .A3(n14758), .A4(n14759), .ZN(
        n14755) );
  NOR4_X1 U9231 ( .A1(n14752), .A2(n14753), .A3(n14754), .A4(n14755), .ZN(
        n14751) );
  NOR2_X1 U9230 ( .A1(n14751), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N139 ) );
  AOI22_X1 U8889 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[31][23] ), .A2(n14249), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[30][23] ), .B2(n17683), .ZN(
        n14408) );
  AOI22_X1 U8888 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[29][23] ), .A2(n17684), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[28][23] ), .B2(n17685), .ZN(
        n14409) );
  AOI222_X1 U8887 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[4][23] ), .A2(n17686), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[25][23] ), .B2(n14245), .C1(
        \pipeline/RegFile_DEC_WB/RegBank[24][23] ), .C2(n17687), .ZN(n14410)
         );
  AOI22_X1 U8886 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[27][23] ), .A2(n14239), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[26][23] ), .B2(n17689), .ZN(
        n14404) );
  AOI22_X1 U8885 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[23][23] ), .A2(n14237), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[22][23] ), .B2(n17691), .ZN(
        n14405) );
  AOI22_X1 U8884 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[21][23] ), .A2(n17692), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[20][23] ), .B2(n17693), .ZN(
        n14406) );
  AOI22_X1 U8883 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[19][23] ), .A2(n17694), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[18][23] ), .B2(n17695), .ZN(
        n14407) );
  NAND4_X1 U8882 ( .A1(n14404), .A2(n14405), .A3(n14406), .A4(n14407), .ZN(
        n14393) );
  AOI22_X1 U8881 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[17][23] ), .A2(n14227), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[16][23] ), .B2(n17697), .ZN(
        n14400) );
  AOI22_X1 U8880 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[12][23] ), .A2(n17698), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[13][23] ), .B2(n17357), .ZN(
        n14401) );
  AOI22_X1 U8879 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[8][23] ), .A2(n17417), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[15][23] ), .B2(n17152), .ZN(
        n14402) );
  AOI22_X1 U8878 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[9][23] ), .A2(n17351), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[10][23] ), .B2(n17699), .ZN(
        n14403) );
  NAND4_X1 U8877 ( .A1(n14400), .A2(n14401), .A3(n14402), .A4(n14403), .ZN(
        n14394) );
  AOI22_X1 U8876 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[11][23] ), .A2(n14215), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[3][23] ), .B2(n17413), .ZN(n14396) );
  AOI22_X1 U8875 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[14][23] ), .A2(n14213), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[5][23] ), .B2(n17414), .ZN(n14397) );
  AOI22_X1 U8874 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[2][23] ), .A2(n17353), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[7][23] ), .B2(n17415), .ZN(n14398) );
  AOI22_X1 U8873 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[6][23] ), .A2(n17354), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[1][23] ), .B2(n17416), .ZN(n14399) );
  NAND4_X1 U8872 ( .A1(n14396), .A2(n14397), .A3(n14398), .A4(n14399), .ZN(
        n14395) );
  NOR4_X1 U8871 ( .A1(n14392), .A2(n14393), .A3(n14394), .A4(n14395), .ZN(
        n14391) );
  NOR2_X1 U8870 ( .A1(n14391), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N157 ) );
  AOI22_X1 U9089 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[31][13] ), .A2(n17154), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[30][13] ), .B2(n17683), .ZN(
        n14608) );
  AOI22_X1 U9088 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[29][13] ), .A2(n17684), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[28][13] ), .B2(n17685), .ZN(
        n14609) );
  AOI222_X1 U9087 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[4][13] ), .A2(n17686), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[25][13] ), .B2(n17153), .C1(
        \pipeline/RegFile_DEC_WB/RegBank[24][13] ), .C2(n17687), .ZN(n14610)
         );
  AOI22_X1 U9086 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[27][13] ), .A2(n17688), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[26][13] ), .B2(n17689), .ZN(
        n14604) );
  AOI22_X1 U9085 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[23][13] ), .A2(n17690), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[22][13] ), .B2(n17691), .ZN(
        n14605) );
  AOI22_X1 U9084 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[21][13] ), .A2(n17692), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[20][13] ), .B2(n17693), .ZN(
        n14606) );
  AOI22_X1 U9083 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[19][13] ), .A2(n17694), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[18][13] ), .B2(n17695), .ZN(
        n14607) );
  NAND4_X1 U9082 ( .A1(n14604), .A2(n14605), .A3(n14606), .A4(n14607), .ZN(
        n14593) );
  AOI22_X1 U9081 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[17][13] ), .A2(n17696), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[16][13] ), .B2(n17697), .ZN(
        n14600) );
  AOI22_X1 U9080 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[12][13] ), .A2(n17698), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[13][13] ), .B2(n14226), .ZN(
        n14601) );
  AOI22_X1 U9079 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[8][13] ), .A2(n14223), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[15][13] ), .B2(n17152), .ZN(
        n14602) );
  AOI22_X1 U9078 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[9][13] ), .A2(n14221), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[10][13] ), .B2(n17699), .ZN(
        n14603) );
  NAND4_X1 U9077 ( .A1(n14600), .A2(n14601), .A3(n14602), .A4(n14603), .ZN(
        n14594) );
  AOI22_X1 U9076 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[11][13] ), .A2(n17151), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[3][13] ), .B2(n14216), .ZN(n14596) );
  AOI22_X1 U9075 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[14][13] ), .A2(n17700), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[5][13] ), .B2(n14214), .ZN(n14597) );
  AOI22_X1 U9074 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[2][13] ), .A2(n17367), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[7][13] ), .B2(n14212), .ZN(n14598) );
  AOI22_X1 U9073 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[6][13] ), .A2(n17368), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[1][13] ), .B2(n14210), .ZN(n14599) );
  NAND4_X1 U9072 ( .A1(n14596), .A2(n14597), .A3(n14598), .A4(n14599), .ZN(
        n14595) );
  NOR4_X1 U9071 ( .A1(n14592), .A2(n14593), .A3(n14594), .A4(n14595), .ZN(
        n14591) );
  NOR2_X1 U9070 ( .A1(n14591), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N147 ) );
  AOI22_X1 U9069 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[31][14] ), .A2(n17154), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[30][14] ), .B2(n17683), .ZN(
        n14588) );
  AOI22_X1 U9068 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[29][14] ), .A2(n17684), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[28][14] ), .B2(n17685), .ZN(
        n14589) );
  AOI222_X1 U9067 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[4][14] ), .A2(n17686), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[25][14] ), .B2(n14245), .C1(
        \pipeline/RegFile_DEC_WB/RegBank[24][14] ), .C2(n17687), .ZN(n14590)
         );
  AOI22_X1 U9066 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[27][14] ), .A2(n17688), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[26][14] ), .B2(n17689), .ZN(
        n14584) );
  AOI22_X1 U9065 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[23][14] ), .A2(n17690), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[22][14] ), .B2(n17691), .ZN(
        n14585) );
  AOI22_X1 U9064 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[21][14] ), .A2(n17692), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[20][14] ), .B2(n17693), .ZN(
        n14586) );
  AOI22_X1 U9063 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[19][14] ), .A2(n17694), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[18][14] ), .B2(n17695), .ZN(
        n14587) );
  NAND4_X1 U9062 ( .A1(n14584), .A2(n14585), .A3(n14586), .A4(n14587), .ZN(
        n14573) );
  AOI22_X1 U9061 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[17][14] ), .A2(n17696), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[16][14] ), .B2(n17697), .ZN(
        n14580) );
  AOI22_X1 U9060 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[12][14] ), .A2(n17698), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[13][14] ), .B2(n17358), .ZN(
        n14581) );
  AOI22_X1 U9059 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[8][14] ), .A2(n14223), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[15][14] ), .B2(n17152), .ZN(
        n14582) );
  AOI22_X1 U9058 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[9][14] ), .A2(n17352), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[10][14] ), .B2(n17699), .ZN(
        n14583) );
  NAND4_X1 U9057 ( .A1(n14580), .A2(n14581), .A3(n14582), .A4(n14583), .ZN(
        n14574) );
  AOI22_X1 U9056 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[11][14] ), .A2(n14215), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[3][14] ), .B2(n14216), .ZN(n14576) );
  AOI22_X1 U9055 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[14][14] ), .A2(n14213), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[5][14] ), .B2(n14214), .ZN(n14577) );
  AOI22_X1 U9054 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[2][14] ), .A2(n17355), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[7][14] ), .B2(n14212), .ZN(n14578) );
  AOI22_X1 U9053 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[6][14] ), .A2(n17356), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[1][14] ), .B2(n14210), .ZN(n14579) );
  NAND4_X1 U9052 ( .A1(n14576), .A2(n14577), .A3(n14578), .A4(n14579), .ZN(
        n14575) );
  NOR4_X1 U9051 ( .A1(n14572), .A2(n14573), .A3(n14574), .A4(n14575), .ZN(
        n14571) );
  NOR2_X1 U9050 ( .A1(n14571), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N148 ) );
  AOI22_X1 U8729 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[31][31] ), .A2(n14249), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[30][31] ), .B2(n14250), .ZN(
        n14241) );
  AOI22_X1 U8728 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[29][31] ), .A2(n14247), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[28][31] ), .B2(n14248), .ZN(
        n14242) );
  AOI222_X1 U8727 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[4][31] ), .A2(n14244), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[25][31] ), .B2(n14245), .C1(
        \pipeline/RegFile_DEC_WB/RegBank[24][31] ), .C2(n17687), .ZN(n14243)
         );
  AOI22_X1 U8726 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[27][31] ), .A2(n14239), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[26][31] ), .B2(n14240), .ZN(
        n14229) );
  AOI22_X1 U8725 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[23][31] ), .A2(n14237), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[22][31] ), .B2(n14238), .ZN(
        n14230) );
  AOI22_X1 U8724 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[21][31] ), .A2(n14235), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[20][31] ), .B2(n14236), .ZN(
        n14231) );
  AOI22_X1 U8723 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[19][31] ), .A2(n14233), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[18][31] ), .B2(n14234), .ZN(
        n14232) );
  NAND4_X1 U8722 ( .A1(n14229), .A2(n14230), .A3(n14231), .A4(n14232), .ZN(
        n14202) );
  AOI22_X1 U8721 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[17][31] ), .A2(n14227), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[16][31] ), .B2(n14228), .ZN(
        n14217) );
  AOI22_X1 U8720 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[12][31] ), .A2(n14225), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[13][31] ), .B2(n17358), .ZN(
        n14218) );
  AOI22_X1 U8719 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[8][31] ), .A2(n14223), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[15][31] ), .B2(n17152), .ZN(
        n14219) );
  AOI22_X1 U8718 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[9][31] ), .A2(n17352), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[10][31] ), .B2(n14222), .ZN(
        n14220) );
  NAND4_X1 U8717 ( .A1(n14217), .A2(n14218), .A3(n14219), .A4(n14220), .ZN(
        n14203) );
  AOI22_X1 U8716 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[11][31] ), .A2(n17151), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[3][31] ), .B2(n14216), .ZN(n14205) );
  AOI22_X1 U8715 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[14][31] ), .A2(n17700), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[5][31] ), .B2(n14214), .ZN(n14206) );
  AOI22_X1 U8714 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[2][31] ), .A2(n17355), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[7][31] ), .B2(n14212), .ZN(n14207) );
  AOI22_X1 U8713 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[6][31] ), .A2(n17356), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[1][31] ), .B2(n14210), .ZN(n14208) );
  NAND4_X1 U8712 ( .A1(n14205), .A2(n14206), .A3(n14207), .A4(n14208), .ZN(
        n14204) );
  NOR4_X1 U8711 ( .A1(n14201), .A2(n14202), .A3(n14203), .A4(n14204), .ZN(
        n14200) );
  NOR2_X1 U8710 ( .A1(n14200), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N165 ) );
  AOI22_X1 U9149 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[31][10] ), .A2(n17154), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[30][10] ), .B2(n17683), .ZN(
        n14668) );
  AOI22_X1 U9148 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[29][10] ), .A2(n17684), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[28][10] ), .B2(n17685), .ZN(
        n14669) );
  AOI222_X1 U9147 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[4][10] ), .A2(n17686), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[25][10] ), .B2(n17153), .C1(
        \pipeline/RegFile_DEC_WB/RegBank[24][10] ), .C2(n17687), .ZN(n14670)
         );
  AOI22_X1 U9146 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[27][10] ), .A2(n17688), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[26][10] ), .B2(n17689), .ZN(
        n14664) );
  AOI22_X1 U9145 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[23][10] ), .A2(n17690), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[22][10] ), .B2(n17691), .ZN(
        n14665) );
  AOI22_X1 U9144 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[21][10] ), .A2(n17692), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[20][10] ), .B2(n17693), .ZN(
        n14666) );
  AOI22_X1 U9143 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[19][10] ), .A2(n17694), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[18][10] ), .B2(n17695), .ZN(
        n14667) );
  NAND4_X1 U9142 ( .A1(n14664), .A2(n14665), .A3(n14666), .A4(n14667), .ZN(
        n14653) );
  AOI22_X1 U9141 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[17][10] ), .A2(n17696), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[16][10] ), .B2(n17697), .ZN(
        n14660) );
  AOI22_X1 U9140 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[12][10] ), .A2(n17698), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[13][10] ), .B2(n17358), .ZN(
        n14661) );
  AOI22_X1 U9139 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[8][10] ), .A2(n14223), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[15][10] ), .B2(n17152), .ZN(
        n14662) );
  AOI22_X1 U9138 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[9][10] ), .A2(n17352), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[10][10] ), .B2(n17699), .ZN(
        n14663) );
  NAND4_X1 U9137 ( .A1(n14660), .A2(n14661), .A3(n14662), .A4(n14663), .ZN(
        n14654) );
  AOI22_X1 U9136 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[11][10] ), .A2(n17151), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[3][10] ), .B2(n14216), .ZN(n14656) );
  AOI22_X1 U9135 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[14][10] ), .A2(n17700), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[5][10] ), .B2(n14214), .ZN(n14657) );
  AOI22_X1 U9134 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[2][10] ), .A2(n17355), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[7][10] ), .B2(n14212), .ZN(n14658) );
  AOI22_X1 U9133 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[6][10] ), .A2(n17356), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[1][10] ), .B2(n14210), .ZN(n14659) );
  NAND4_X1 U9132 ( .A1(n14656), .A2(n14657), .A3(n14658), .A4(n14659), .ZN(
        n14655) );
  NOR4_X1 U9131 ( .A1(n14652), .A2(n14653), .A3(n14654), .A4(n14655), .ZN(
        n14651) );
  NOR2_X1 U9130 ( .A1(n14651), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N144 ) );
  AOI22_X1 U8829 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[31][26] ), .A2(n17154), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[30][26] ), .B2(n17683), .ZN(
        n14348) );
  AOI22_X1 U8828 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[29][26] ), .A2(n17684), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[28][26] ), .B2(n17685), .ZN(
        n14349) );
  AOI222_X1 U8827 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[4][26] ), .A2(n17686), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[25][26] ), .B2(n17153), .C1(
        \pipeline/RegFile_DEC_WB/RegBank[24][26] ), .C2(n17687), .ZN(n14350)
         );
  AOI22_X1 U8826 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[27][26] ), .A2(n17688), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[26][26] ), .B2(n17689), .ZN(
        n14344) );
  AOI22_X1 U8825 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[23][26] ), .A2(n17690), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[22][26] ), .B2(n17691), .ZN(
        n14345) );
  AOI22_X1 U8824 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[21][26] ), .A2(n17692), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[20][26] ), .B2(n17693), .ZN(
        n14346) );
  AOI22_X1 U8823 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[19][26] ), .A2(n17694), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[18][26] ), .B2(n17695), .ZN(
        n14347) );
  NAND4_X1 U8822 ( .A1(n14344), .A2(n14345), .A3(n14346), .A4(n14347), .ZN(
        n14333) );
  AOI22_X1 U8821 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[17][26] ), .A2(n17696), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[16][26] ), .B2(n17697), .ZN(
        n14340) );
  AOI22_X1 U8820 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[12][26] ), .A2(n17698), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[13][26] ), .B2(n17357), .ZN(
        n14341) );
  AOI22_X1 U8819 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[8][26] ), .A2(n17417), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[15][26] ), .B2(n14224), .ZN(
        n14342) );
  AOI22_X1 U8818 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[9][26] ), .A2(n17351), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[10][26] ), .B2(n17699), .ZN(
        n14343) );
  NAND4_X1 U8817 ( .A1(n14340), .A2(n14341), .A3(n14342), .A4(n14343), .ZN(
        n14334) );
  AOI22_X1 U8816 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[11][26] ), .A2(n17151), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[3][26] ), .B2(n17413), .ZN(n14336) );
  AOI22_X1 U8815 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[14][26] ), .A2(n17700), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[5][26] ), .B2(n17414), .ZN(n14337) );
  AOI22_X1 U8814 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[2][26] ), .A2(n17353), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[7][26] ), .B2(n17415), .ZN(n14338) );
  AOI22_X1 U8813 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[6][26] ), .A2(n17354), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[1][26] ), .B2(n17416), .ZN(n14339) );
  NAND4_X1 U8812 ( .A1(n14336), .A2(n14337), .A3(n14338), .A4(n14339), .ZN(
        n14335) );
  NOR4_X1 U8811 ( .A1(n14332), .A2(n14333), .A3(n14334), .A4(n14335), .ZN(
        n14331) );
  NOR2_X1 U8810 ( .A1(n14331), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N160 ) );
  AOI22_X1 U9329 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[31][1] ), .A2(n17154), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[30][1] ), .B2(n17683), .ZN(n14848) );
  AOI22_X1 U9328 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[29][1] ), .A2(n17684), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[28][1] ), .B2(n17685), .ZN(n14849) );
  AOI222_X1 U9327 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[4][1] ), .A2(n17686), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[25][1] ), .B2(n17153), .C1(
        \pipeline/RegFile_DEC_WB/RegBank[24][1] ), .C2(n17687), .ZN(n14850) );
  AOI22_X1 U9326 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[27][1] ), .A2(n17688), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[26][1] ), .B2(n17689), .ZN(n14844) );
  AOI22_X1 U9325 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[23][1] ), .A2(n17690), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[22][1] ), .B2(n17691), .ZN(n14845) );
  AOI22_X1 U9324 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[21][1] ), .A2(n17692), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[20][1] ), .B2(n17693), .ZN(n14846) );
  AOI22_X1 U9323 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[19][1] ), .A2(n17694), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[18][1] ), .B2(n17695), .ZN(n14847) );
  NAND4_X1 U9322 ( .A1(n14844), .A2(n14845), .A3(n14846), .A4(n14847), .ZN(
        n14833) );
  AOI22_X1 U9321 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[17][1] ), .A2(n17696), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[16][1] ), .B2(n17697), .ZN(n14840) );
  AOI22_X1 U9320 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[12][1] ), .A2(n17698), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[13][1] ), .B2(n17357), .ZN(n14841) );
  AOI22_X1 U9319 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[8][1] ), .A2(n17417), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[15][1] ), .B2(n14224), .ZN(n14842) );
  AOI22_X1 U9318 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[9][1] ), .A2(n17351), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[10][1] ), .B2(n17699), .ZN(n14843) );
  NAND4_X1 U9317 ( .A1(n14840), .A2(n14841), .A3(n14842), .A4(n14843), .ZN(
        n14834) );
  AOI22_X1 U9316 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[11][1] ), .A2(n17151), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[3][1] ), .B2(n17413), .ZN(n14836)
         );
  AOI22_X1 U9315 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[14][1] ), .A2(n17700), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[5][1] ), .B2(n17414), .ZN(n14837)
         );
  AOI22_X1 U9314 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[2][1] ), .A2(n17353), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[7][1] ), .B2(n17415), .ZN(n14838)
         );
  AOI22_X1 U9313 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[6][1] ), .A2(n17354), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[1][1] ), .B2(n17416), .ZN(n14839)
         );
  NAND4_X1 U9312 ( .A1(n14836), .A2(n14837), .A3(n14838), .A4(n14839), .ZN(
        n14835) );
  NOR4_X1 U9311 ( .A1(n14832), .A2(n14833), .A3(n14834), .A4(n14835), .ZN(
        n14831) );
  NOR2_X1 U9310 ( .A1(n14831), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N135 ) );
  AOI22_X1 U8789 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[31][28] ), .A2(n17154), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[30][28] ), .B2(n17683), .ZN(
        n14308) );
  AOI22_X1 U8788 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[29][28] ), .A2(n17684), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[28][28] ), .B2(n17685), .ZN(
        n14309) );
  AOI222_X1 U8787 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[4][28] ), .A2(n17686), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[25][28] ), .B2(n17153), .C1(
        \pipeline/RegFile_DEC_WB/RegBank[24][28] ), .C2(n17687), .ZN(n14310)
         );
  AOI22_X1 U8786 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[27][28] ), .A2(n17688), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[26][28] ), .B2(n17689), .ZN(
        n14304) );
  AOI22_X1 U8785 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[23][28] ), .A2(n17690), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[22][28] ), .B2(n17691), .ZN(
        n14305) );
  AOI22_X1 U8784 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[21][28] ), .A2(n17692), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[20][28] ), .B2(n17693), .ZN(
        n14306) );
  AOI22_X1 U8783 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[19][28] ), .A2(n17694), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[18][28] ), .B2(n17695), .ZN(
        n14307) );
  NAND4_X1 U8782 ( .A1(n14304), .A2(n14305), .A3(n14306), .A4(n14307), .ZN(
        n14293) );
  AOI22_X1 U8781 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[17][28] ), .A2(n17696), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[16][28] ), .B2(n17697), .ZN(
        n14300) );
  AOI22_X1 U8780 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[12][28] ), .A2(n17698), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[13][28] ), .B2(n17358), .ZN(
        n14301) );
  AOI22_X1 U8779 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[8][28] ), .A2(n17417), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[15][28] ), .B2(n14224), .ZN(
        n14302) );
  AOI22_X1 U8778 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[9][28] ), .A2(n17352), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[10][28] ), .B2(n17699), .ZN(
        n14303) );
  NAND4_X1 U8777 ( .A1(n14300), .A2(n14301), .A3(n14302), .A4(n14303), .ZN(
        n14294) );
  AOI22_X1 U8776 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[11][28] ), .A2(n17151), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[3][28] ), .B2(n17413), .ZN(n14296) );
  AOI22_X1 U8775 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[14][28] ), .A2(n17700), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[5][28] ), .B2(n17414), .ZN(n14297) );
  AOI22_X1 U8774 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[2][28] ), .A2(n17355), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[7][28] ), .B2(n17415), .ZN(n14298) );
  AOI22_X1 U8773 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[6][28] ), .A2(n17356), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[1][28] ), .B2(n17416), .ZN(n14299) );
  NAND4_X1 U8772 ( .A1(n14296), .A2(n14297), .A3(n14298), .A4(n14299), .ZN(
        n14295) );
  NOR4_X1 U8771 ( .A1(n14292), .A2(n14293), .A3(n14294), .A4(n14295), .ZN(
        n14291) );
  NOR2_X1 U8770 ( .A1(n14291), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N162 ) );
  AOI22_X1 U9189 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[31][8] ), .A2(n17154), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[30][8] ), .B2(n17683), .ZN(n14708) );
  AOI22_X1 U9188 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[29][8] ), .A2(n17684), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[28][8] ), .B2(n17685), .ZN(n14709) );
  AOI222_X1 U9187 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[4][8] ), .A2(n17686), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[25][8] ), .B2(n17153), .C1(
        \pipeline/RegFile_DEC_WB/RegBank[24][8] ), .C2(n17687), .ZN(n14710) );
  AOI22_X1 U9186 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[27][8] ), .A2(n17688), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[26][8] ), .B2(n17689), .ZN(n14704) );
  AOI22_X1 U9185 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[23][8] ), .A2(n17690), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[22][8] ), .B2(n17691), .ZN(n14705) );
  AOI22_X1 U9184 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[21][8] ), .A2(n17692), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[20][8] ), .B2(n17693), .ZN(n14706) );
  AOI22_X1 U9183 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[19][8] ), .A2(n17694), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[18][8] ), .B2(n17695), .ZN(n14707) );
  NAND4_X1 U9182 ( .A1(n14704), .A2(n14705), .A3(n14706), .A4(n14707), .ZN(
        n14693) );
  AOI22_X1 U9181 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[17][8] ), .A2(n17696), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[16][8] ), .B2(n17697), .ZN(n14700) );
  AOI22_X1 U9180 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[12][8] ), .A2(n17698), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[13][8] ), .B2(n17358), .ZN(n14701) );
  AOI22_X1 U9179 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[8][8] ), .A2(n17417), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[15][8] ), .B2(n17152), .ZN(n14702) );
  AOI22_X1 U9178 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[9][8] ), .A2(n17352), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[10][8] ), .B2(n17699), .ZN(n14703) );
  NAND4_X1 U9177 ( .A1(n14700), .A2(n14701), .A3(n14702), .A4(n14703), .ZN(
        n14694) );
  AOI22_X1 U9176 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[11][8] ), .A2(n17151), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[3][8] ), .B2(n17413), .ZN(n14696)
         );
  AOI22_X1 U9175 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[14][8] ), .A2(n17700), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[5][8] ), .B2(n17414), .ZN(n14697)
         );
  AOI22_X1 U9174 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[2][8] ), .A2(n17355), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[7][8] ), .B2(n17415), .ZN(n14698)
         );
  AOI22_X1 U9173 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[6][8] ), .A2(n17356), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[1][8] ), .B2(n17416), .ZN(n14699)
         );
  NAND4_X1 U9172 ( .A1(n14696), .A2(n14697), .A3(n14698), .A4(n14699), .ZN(
        n14695) );
  NOR4_X1 U9171 ( .A1(n14692), .A2(n14693), .A3(n14694), .A4(n14695), .ZN(
        n14691) );
  NOR2_X1 U9170 ( .A1(n14691), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N142 ) );
  AOI22_X1 U8869 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[31][24] ), .A2(n17154), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[30][24] ), .B2(n17683), .ZN(
        n14388) );
  AOI22_X1 U8868 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[29][24] ), .A2(n17684), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[28][24] ), .B2(n17685), .ZN(
        n14389) );
  AOI222_X1 U8867 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[4][24] ), .A2(n17686), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[25][24] ), .B2(n17153), .C1(
        \pipeline/RegFile_DEC_WB/RegBank[24][24] ), .C2(n17687), .ZN(n14390)
         );
  AOI22_X1 U8866 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[27][24] ), .A2(n17688), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[26][24] ), .B2(n17689), .ZN(
        n14384) );
  AOI22_X1 U8865 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[23][24] ), .A2(n17690), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[22][24] ), .B2(n17691), .ZN(
        n14385) );
  AOI22_X1 U8864 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[21][24] ), .A2(n17692), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[20][24] ), .B2(n17693), .ZN(
        n14386) );
  AOI22_X1 U8863 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[19][24] ), .A2(n17694), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[18][24] ), .B2(n17695), .ZN(
        n14387) );
  NAND4_X1 U8862 ( .A1(n14384), .A2(n14385), .A3(n14386), .A4(n14387), .ZN(
        n14373) );
  AOI22_X1 U8861 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[17][24] ), .A2(n17696), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[16][24] ), .B2(n17697), .ZN(
        n14380) );
  AOI22_X1 U8860 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[12][24] ), .A2(n17698), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[13][24] ), .B2(n17357), .ZN(
        n14381) );
  AOI22_X1 U8859 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[8][24] ), .A2(n17417), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[15][24] ), .B2(n14224), .ZN(
        n14382) );
  AOI22_X1 U8858 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[9][24] ), .A2(n17351), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[10][24] ), .B2(n17699), .ZN(
        n14383) );
  NAND4_X1 U8857 ( .A1(n14380), .A2(n14381), .A3(n14382), .A4(n14383), .ZN(
        n14374) );
  AOI22_X1 U8856 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[11][24] ), .A2(n17151), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[3][24] ), .B2(n17413), .ZN(n14376) );
  AOI22_X1 U8855 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[14][24] ), .A2(n17700), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[5][24] ), .B2(n17414), .ZN(n14377) );
  AOI22_X1 U8854 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[2][24] ), .A2(n17353), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[7][24] ), .B2(n17415), .ZN(n14378) );
  AOI22_X1 U8853 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[6][24] ), .A2(n17354), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[1][24] ), .B2(n17416), .ZN(n14379) );
  NAND4_X1 U8852 ( .A1(n14376), .A2(n14377), .A3(n14378), .A4(n14379), .ZN(
        n14375) );
  NOR4_X1 U8851 ( .A1(n14372), .A2(n14373), .A3(n14374), .A4(n14375), .ZN(
        n14371) );
  NOR2_X1 U8850 ( .A1(n14371), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N158 ) );
  AOI22_X1 U9309 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[31][2] ), .A2(n17154), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[30][2] ), .B2(n17683), .ZN(n14828) );
  AOI22_X1 U9308 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[29][2] ), .A2(n17684), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[28][2] ), .B2(n17685), .ZN(n14829) );
  AOI222_X1 U9307 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[4][2] ), .A2(n14244), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[25][2] ), .B2(n17153), .C1(
        \pipeline/RegFile_DEC_WB/RegBank[24][2] ), .C2(n14246), .ZN(n14830) );
  AOI22_X1 U9306 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[27][2] ), .A2(n17688), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[26][2] ), .B2(n14240), .ZN(n14824) );
  AOI22_X1 U9305 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[23][2] ), .A2(n17690), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[22][2] ), .B2(n17691), .ZN(n14825) );
  AOI22_X1 U9304 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[21][2] ), .A2(n17692), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[20][2] ), .B2(n14236), .ZN(n14826) );
  AOI22_X1 U9303 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[19][2] ), .A2(n17694), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[18][2] ), .B2(n17695), .ZN(n14827) );
  NAND4_X1 U9302 ( .A1(n14824), .A2(n14825), .A3(n14826), .A4(n14827), .ZN(
        n14813) );
  AOI22_X1 U9301 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[17][2] ), .A2(n17696), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[16][2] ), .B2(n14228), .ZN(n14820) );
  AOI22_X1 U9300 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[12][2] ), .A2(n17698), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[13][2] ), .B2(n17357), .ZN(n14821) );
  AOI22_X1 U9299 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[8][2] ), .A2(n17417), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[15][2] ), .B2(n17152), .ZN(n14822) );
  AOI22_X1 U9298 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[9][2] ), .A2(n17351), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[10][2] ), .B2(n17699), .ZN(n14823) );
  NAND4_X1 U9297 ( .A1(n14820), .A2(n14821), .A3(n14822), .A4(n14823), .ZN(
        n14814) );
  AOI22_X1 U9296 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[11][2] ), .A2(n17151), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[3][2] ), .B2(n17413), .ZN(n14816)
         );
  AOI22_X1 U9295 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[14][2] ), .A2(n17700), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[5][2] ), .B2(n17414), .ZN(n14817)
         );
  AOI22_X1 U9294 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[2][2] ), .A2(n17353), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[7][2] ), .B2(n17415), .ZN(n14818)
         );
  AOI22_X1 U9293 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[6][2] ), .A2(n17354), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[1][2] ), .B2(n17416), .ZN(n14819)
         );
  NAND4_X1 U9292 ( .A1(n14816), .A2(n14817), .A3(n14818), .A4(n14819), .ZN(
        n14815) );
  NOR4_X1 U9291 ( .A1(n14812), .A2(n14813), .A3(n14814), .A4(n14815), .ZN(
        n14811) );
  AOI21_X1 U9290 ( .B1(n14025), .B2(n14811), .A(n14168), .ZN(
        \pipeline/IDEX_Stage/N136 ) );
  NOR2_X1 U8655 ( .A1(n17313), .A2(n14059), .ZN(n14084) );
  NAND2_X1 U8653 ( .A1(\pipeline/inst_IFID_DEC[29] ), .A2(n14190), .ZN(n13998)
         );
  NOR2_X1 U8651 ( .A1(n17347), .A2(n14058), .ZN(n13999) );
  NAND2_X1 U8650 ( .A1(\pipeline/inst_IFID_DEC[30] ), .A2(
        \pipeline/inst_IFID_DEC[26] ), .ZN(n14189) );
  NOR4_X1 U8649 ( .A1(\pipeline/inst_IFID_DEC[27] ), .A2(n17382), .A3(n17348), 
        .A4(n14189), .ZN(n14040) );
  NOR2_X1 U8648 ( .A1(n13999), .A2(n14040), .ZN(n14042) );
  NAND2_X1 U8647 ( .A1(n17313), .A2(n14001), .ZN(n14011) );
  NAND2_X1 U8645 ( .A1(\pipeline/inst_IFID_DEC[30] ), .A2(n14185), .ZN(n13997)
         );
  NAND2_X1 U8644 ( .A1(n14042), .A2(n13997), .ZN(n14016) );
  NOR4_X1 U8643 ( .A1(n17313), .A2(n17347), .A3(n17382), .A4(
        \pipeline/inst_IFID_DEC[28] ), .ZN(n14022) );
  NOR2_X1 U8642 ( .A1(n14016), .A2(n14022), .ZN(n14188) );
  NAND2_X1 U8641 ( .A1(n14029), .A2(n14188), .ZN(n14009) );
  NAND2_X1 U8640 ( .A1(n14049), .A2(\pipeline/inst_IFID_DEC[29] ), .ZN(n14187)
         );
  AOI21_X1 U8639 ( .B1(\pipeline/inst_IFID_DEC[27] ), .B2(n14176), .A(n14187), 
        .ZN(n14183) );
  NAND2_X1 U8638 ( .A1(\pipeline/inst_IFID_DEC[30] ), .A2(n17409), .ZN(n14047)
         );
  NOR2_X1 U8637 ( .A1(n14186), .A2(n14047), .ZN(n14061) );
  AOI21_X1 U8636 ( .B1(n14185), .B2(n17347), .A(n14061), .ZN(n14028) );
  NAND4_X1 U8635 ( .A1(n14049), .A2(n17382), .A3(\pipeline/inst_IFID_DEC[27] ), 
        .A4(\pipeline/inst_IFID_DEC[30] ), .ZN(n14019) );
  NAND2_X1 U8634 ( .A1(n14028), .A2(n14019), .ZN(n14184) );
  NAND2_X1 U8632 ( .A1(\pipeline/stageD/offset_to_jump_temp [5]), .A2(n17404), 
        .ZN(n14181) );
  NOR3_X1 U8631 ( .A1(\pipeline/stageD/offset_to_jump_temp [4]), .A2(
        \pipeline/stageD/offset_to_jump_temp [3]), .A3(n17404), .ZN(n14067) );
  NAND2_X1 U8628 ( .A1(n14179), .A2(n14051), .ZN(n14024) );
  OAI211_X1 U8627 ( .C1(\pipeline/stageD/offset_to_jump_temp [4]), .C2(n14181), 
        .A(n14066), .B(n14024), .ZN(n14172) );
  NOR2_X1 U8625 ( .A1(n17406), .A2(n17076), .ZN(n14031) );
  OAI221_X1 U8624 ( .B1(n14032), .B2(n14031), .C1(n14032), .C2(n17350), .A(
        n14067), .ZN(n14178) );
  NOR2_X1 U8621 ( .A1(\pipeline/stageD/offset_to_jump_temp [4]), .A2(n14180), 
        .ZN(n14065) );
  NOR2_X1 U8619 ( .A1(n17076), .A2(n14180), .ZN(n14045) );
  AOI21_X1 U8618 ( .B1(n14031), .B2(n14179), .A(n14045), .ZN(n14023) );
  NAND2_X1 U8617 ( .A1(n14051), .A2(n14067), .ZN(n14064) );
  NAND4_X1 U8616 ( .A1(n14178), .A2(n14006), .A3(n14023), .A4(n14064), .ZN(
        n14173) );
  OAI21_X1 U8613 ( .B1(n14172), .B2(n14173), .A(n14005), .ZN(n14170) );
  OAI221_X1 U8612 ( .B1(n14168), .B2(n13980), .C1(n14168), .C2(n14170), .A(
        n17682), .ZN(\pipeline/IDEX_Stage/N90 ) );
  OAI22_X1 U9438 ( .A1(n14931), .A2(n17075), .B1(n17109), .B2(n17468), .ZN(
        \pipeline/IDEX_Stage/N109 ) );
  OAI22_X1 U9430 ( .A1(n14923), .A2(n17075), .B1(n17682), .B2(n17441), .ZN(
        \pipeline/IDEX_Stage/N113 ) );
  OAI22_X1 U9412 ( .A1(n14905), .A2(n17075), .B1(n17682), .B2(n17463), .ZN(
        \pipeline/IDEX_Stage/N122 ) );
  OAI22_X1 U9446 ( .A1(n14939), .A2(n17075), .B1(n17109), .B2(n17439), .ZN(
        \pipeline/IDEX_Stage/N105 ) );
  OAI22_X1 U9428 ( .A1(n14921), .A2(n17075), .B1(n17109), .B2(n17459), .ZN(
        \pipeline/IDEX_Stage/N114 ) );
  OAI22_X1 U9436 ( .A1(n14929), .A2(n17075), .B1(n17109), .B2(n17457), .ZN(
        \pipeline/IDEX_Stage/N110 ) );
  OAI22_X1 U9410 ( .A1(n14903), .A2(n17075), .B1(n17109), .B2(n17448), .ZN(
        \pipeline/IDEX_Stage/N123 ) );
  OAI22_X1 U9418 ( .A1(n14911), .A2(n17075), .B1(n17109), .B2(n17443), .ZN(
        \pipeline/IDEX_Stage/N119 ) );
  OAI22_X1 U9444 ( .A1(n14937), .A2(n17075), .B1(n17109), .B2(n17455), .ZN(
        \pipeline/IDEX_Stage/N106 ) );
  OAI22_X1 U9400 ( .A1(n14893), .A2(n17075), .B1(n17682), .B2(n17466), .ZN(
        \pipeline/IDEX_Stage/N128 ) );
  OAI22_X1 U9440 ( .A1(n14933), .A2(n17075), .B1(n17682), .B2(n17456), .ZN(
        \pipeline/IDEX_Stage/N108 ) );
  OAI22_X1 U9398 ( .A1(n14891), .A2(n17075), .B1(n17682), .B2(n17469), .ZN(
        \pipeline/IDEX_Stage/N129 ) );
  OAI22_X1 U9450 ( .A1(n14943), .A2(n17075), .B1(n17109), .B2(n17446), .ZN(
        \pipeline/IDEX_Stage/N103 ) );
  OAI22_X1 U9406 ( .A1(n14899), .A2(n17075), .B1(n17682), .B2(n17435), .ZN(
        \pipeline/IDEX_Stage/N125 ) );
  OAI22_X1 U9404 ( .A1(n14897), .A2(n17075), .B1(n17682), .B2(n17465), .ZN(
        \pipeline/IDEX_Stage/N126 ) );
  OAI22_X1 U9448 ( .A1(n14941), .A2(n17075), .B1(n17682), .B2(n17470), .ZN(
        \pipeline/IDEX_Stage/N104 ) );
  OAI22_X1 U9396 ( .A1(n14889), .A2(n17075), .B1(n17109), .B2(n17467), .ZN(
        \pipeline/IDEX_Stage/N130 ) );
  OAI22_X1 U9434 ( .A1(n14927), .A2(n17075), .B1(n17109), .B2(n17436), .ZN(
        \pipeline/IDEX_Stage/N111 ) );
  OAI22_X1 U9426 ( .A1(n14919), .A2(n17075), .B1(n17109), .B2(n17442), .ZN(
        \pipeline/IDEX_Stage/N115 ) );
  OAI22_X1 U9392 ( .A1(n14885), .A2(n17075), .B1(n17109), .B2(n17471), .ZN(
        \pipeline/IDEX_Stage/N132 ) );
  OAI22_X1 U9432 ( .A1(n14925), .A2(n17075), .B1(n17109), .B2(n17458), .ZN(
        \pipeline/IDEX_Stage/N112 ) );
  OAI22_X1 U9416 ( .A1(n14909), .A2(n17075), .B1(n17109), .B2(n17462), .ZN(
        \pipeline/IDEX_Stage/N120 ) );
  OAI22_X1 U9408 ( .A1(n14901), .A2(n17075), .B1(n17109), .B2(n17464), .ZN(
        \pipeline/IDEX_Stage/N124 ) );
  AOI22_X1 U8949 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[31][20] ), .A2(n17154), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[30][20] ), .B2(n17683), .ZN(
        n14468) );
  AOI22_X1 U8948 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[29][20] ), .A2(n17684), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[28][20] ), .B2(n17685), .ZN(
        n14469) );
  AOI222_X1 U8947 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[4][20] ), .A2(n14244), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[25][20] ), .B2(n17153), .C1(
        \pipeline/RegFile_DEC_WB/RegBank[24][20] ), .C2(n14246), .ZN(n14470)
         );
  AOI22_X1 U8946 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[27][20] ), .A2(n17688), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[26][20] ), .B2(n14240), .ZN(
        n14464) );
  AOI22_X1 U8945 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[23][20] ), .A2(n17690), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[22][20] ), .B2(n17691), .ZN(
        n14465) );
  AOI22_X1 U8944 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[21][20] ), .A2(n17692), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[20][20] ), .B2(n14236), .ZN(
        n14466) );
  AOI22_X1 U8943 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[19][20] ), .A2(n17694), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[18][20] ), .B2(n17695), .ZN(
        n14467) );
  NAND4_X1 U8942 ( .A1(n14464), .A2(n14465), .A3(n14466), .A4(n14467), .ZN(
        n14453) );
  AOI22_X1 U8941 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[17][20] ), .A2(n17696), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[16][20] ), .B2(n14228), .ZN(
        n14460) );
  AOI22_X1 U8940 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[12][20] ), .A2(n17698), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[13][20] ), .B2(n14226), .ZN(
        n14461) );
  AOI22_X1 U8939 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[8][20] ), .A2(n14223), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[15][20] ), .B2(n17152), .ZN(
        n14462) );
  AOI22_X1 U8938 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[9][20] ), .A2(n14221), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[10][20] ), .B2(n17699), .ZN(
        n14463) );
  NAND4_X1 U8937 ( .A1(n14460), .A2(n14461), .A3(n14462), .A4(n14463), .ZN(
        n14454) );
  AOI22_X1 U8936 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[11][20] ), .A2(n17151), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[3][20] ), .B2(n14216), .ZN(n14456) );
  AOI22_X1 U8935 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[14][20] ), .A2(n17700), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[5][20] ), .B2(n14214), .ZN(n14457) );
  AOI22_X1 U8934 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[2][20] ), .A2(n17367), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[7][20] ), .B2(n14212), .ZN(n14458) );
  AOI22_X1 U8933 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[6][20] ), .A2(n17368), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[1][20] ), .B2(n14210), .ZN(n14459) );
  NAND4_X1 U8932 ( .A1(n14456), .A2(n14457), .A3(n14458), .A4(n14459), .ZN(
        n14455) );
  NOR4_X1 U8931 ( .A1(n14452), .A2(n14453), .A3(n14454), .A4(n14455), .ZN(
        n14451) );
  NOR2_X1 U8930 ( .A1(n14451), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N154 ) );
  AOI22_X1 U8929 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[31][21] ), .A2(n17154), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[30][21] ), .B2(n14250), .ZN(
        n14448) );
  AOI22_X1 U8928 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[29][21] ), .A2(n17684), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[28][21] ), .B2(n14248), .ZN(
        n14449) );
  AOI222_X1 U8927 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[4][21] ), .A2(n17686), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[25][21] ), .B2(n17153), .C1(
        \pipeline/RegFile_DEC_WB/RegBank[24][21] ), .C2(n17687), .ZN(n14450)
         );
  AOI22_X1 U8926 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[27][21] ), .A2(n17688), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[26][21] ), .B2(n17689), .ZN(
        n14444) );
  AOI22_X1 U8925 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[23][21] ), .A2(n17690), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[22][21] ), .B2(n14238), .ZN(
        n14445) );
  AOI22_X1 U8924 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[21][21] ), .A2(n14235), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[20][21] ), .B2(n17693), .ZN(
        n14446) );
  AOI22_X1 U8923 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[19][21] ), .A2(n14233), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[18][21] ), .B2(n17695), .ZN(
        n14447) );
  NAND4_X1 U8922 ( .A1(n14444), .A2(n14445), .A3(n14446), .A4(n14447), .ZN(
        n14433) );
  AOI22_X1 U8921 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[17][21] ), .A2(n17696), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[16][21] ), .B2(n17697), .ZN(
        n14440) );
  AOI22_X1 U8920 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[12][21] ), .A2(n14225), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[13][21] ), .B2(n14226), .ZN(
        n14441) );
  AOI22_X1 U8919 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[8][21] ), .A2(n14223), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[15][21] ), .B2(n17152), .ZN(
        n14442) );
  AOI22_X1 U8918 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[9][21] ), .A2(n14221), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[10][21] ), .B2(n17699), .ZN(
        n14443) );
  NAND4_X1 U8917 ( .A1(n14440), .A2(n14441), .A3(n14442), .A4(n14443), .ZN(
        n14434) );
  AOI22_X1 U8916 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[11][21] ), .A2(n17151), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[3][21] ), .B2(n14216), .ZN(n14436) );
  AOI22_X1 U8915 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[14][21] ), .A2(n14213), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[5][21] ), .B2(n14214), .ZN(n14437) );
  AOI22_X1 U8914 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[2][21] ), .A2(n17367), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[7][21] ), .B2(n14212), .ZN(n14438) );
  AOI22_X1 U8913 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[6][21] ), .A2(n17368), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[1][21] ), .B2(n14210), .ZN(n14439) );
  NAND4_X1 U8912 ( .A1(n14436), .A2(n14437), .A3(n14438), .A4(n14439), .ZN(
        n14435) );
  NOR4_X1 U8911 ( .A1(n14432), .A2(n14433), .A3(n14434), .A4(n14435), .ZN(
        n14431) );
  NOR2_X1 U8910 ( .A1(n14431), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N155 ) );
  AOI22_X1 U9029 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[31][16] ), .A2(n17154), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[30][16] ), .B2(n14250), .ZN(
        n14548) );
  AOI22_X1 U9028 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[29][16] ), .A2(n17684), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[28][16] ), .B2(n14248), .ZN(
        n14549) );
  AOI222_X1 U9027 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[4][16] ), .A2(n14244), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[25][16] ), .B2(n17153), .C1(
        \pipeline/RegFile_DEC_WB/RegBank[24][16] ), .C2(n17687), .ZN(n14550)
         );
  AOI22_X1 U9026 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[27][16] ), .A2(n17688), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[26][16] ), .B2(n14240), .ZN(
        n14544) );
  AOI22_X1 U9025 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[23][16] ), .A2(n17690), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[22][16] ), .B2(n14238), .ZN(
        n14545) );
  AOI22_X1 U9024 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[21][16] ), .A2(n17692), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[20][16] ), .B2(n14236), .ZN(
        n14546) );
  AOI22_X1 U9023 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[19][16] ), .A2(n17694), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[18][16] ), .B2(n14234), .ZN(
        n14547) );
  NAND4_X1 U9022 ( .A1(n14544), .A2(n14545), .A3(n14546), .A4(n14547), .ZN(
        n14533) );
  AOI22_X1 U9021 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[17][16] ), .A2(n17696), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[16][16] ), .B2(n14228), .ZN(
        n14540) );
  AOI22_X1 U9020 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[12][16] ), .A2(n14225), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[13][16] ), .B2(n14226), .ZN(
        n14541) );
  AOI22_X1 U9019 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[8][16] ), .A2(n14223), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[15][16] ), .B2(n17152), .ZN(
        n14542) );
  AOI22_X1 U9018 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[9][16] ), .A2(n14221), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[10][16] ), .B2(n14222), .ZN(
        n14543) );
  NAND4_X1 U9017 ( .A1(n14540), .A2(n14541), .A3(n14542), .A4(n14543), .ZN(
        n14534) );
  AOI22_X1 U9016 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[11][16] ), .A2(n17151), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[3][16] ), .B2(n14216), .ZN(n14536) );
  AOI22_X1 U9015 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[14][16] ), .A2(n14213), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[5][16] ), .B2(n14214), .ZN(n14537) );
  AOI22_X1 U9014 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[2][16] ), .A2(n17367), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[7][16] ), .B2(n14212), .ZN(n14538) );
  AOI22_X1 U9013 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[6][16] ), .A2(n17368), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[1][16] ), .B2(n14210), .ZN(n14539) );
  NAND4_X1 U9012 ( .A1(n14536), .A2(n14537), .A3(n14538), .A4(n14539), .ZN(
        n14535) );
  NOR4_X1 U9011 ( .A1(n14532), .A2(n14533), .A3(n14534), .A4(n14535), .ZN(
        n14531) );
  NOR2_X1 U9010 ( .A1(n14531), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N150 ) );
  AOI22_X1 U9109 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[31][12] ), .A2(n17154), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[30][12] ), .B2(n14250), .ZN(
        n14628) );
  AOI22_X1 U9108 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[29][12] ), .A2(n17684), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[28][12] ), .B2(n14248), .ZN(
        n14629) );
  AOI222_X1 U9107 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[4][12] ), .A2(n17686), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[25][12] ), .B2(n17153), .C1(
        \pipeline/RegFile_DEC_WB/RegBank[24][12] ), .C2(n14246), .ZN(n14630)
         );
  AOI22_X1 U9106 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[27][12] ), .A2(n14239), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[26][12] ), .B2(n17689), .ZN(
        n14624) );
  AOI22_X1 U9105 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[23][12] ), .A2(n17690), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[22][12] ), .B2(n14238), .ZN(
        n14625) );
  AOI22_X1 U9104 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[21][12] ), .A2(n17692), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[20][12] ), .B2(n17693), .ZN(
        n14626) );
  AOI22_X1 U9103 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[19][12] ), .A2(n17694), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[18][12] ), .B2(n14234), .ZN(
        n14627) );
  NAND4_X1 U9102 ( .A1(n14624), .A2(n14625), .A3(n14626), .A4(n14627), .ZN(
        n14613) );
  AOI22_X1 U9101 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[17][12] ), .A2(n14227), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[16][12] ), .B2(n17697), .ZN(
        n14620) );
  AOI22_X1 U9100 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[12][12] ), .A2(n17698), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[13][12] ), .B2(n14226), .ZN(
        n14621) );
  AOI22_X1 U9099 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[8][12] ), .A2(n14223), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[15][12] ), .B2(n17152), .ZN(
        n14622) );
  AOI22_X1 U9098 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[9][12] ), .A2(n14221), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[10][12] ), .B2(n14222), .ZN(
        n14623) );
  NAND4_X1 U9097 ( .A1(n14620), .A2(n14621), .A3(n14622), .A4(n14623), .ZN(
        n14614) );
  AOI22_X1 U9096 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[11][12] ), .A2(n17151), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[3][12] ), .B2(n14216), .ZN(n14616) );
  AOI22_X1 U9095 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[14][12] ), .A2(n14213), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[5][12] ), .B2(n14214), .ZN(n14617) );
  AOI22_X1 U9094 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[2][12] ), .A2(n17367), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[7][12] ), .B2(n14212), .ZN(n14618) );
  AOI22_X1 U9093 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[6][12] ), .A2(n17368), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[1][12] ), .B2(n14210), .ZN(n14619) );
  NAND4_X1 U9092 ( .A1(n14616), .A2(n14617), .A3(n14618), .A4(n14619), .ZN(
        n14615) );
  NOR4_X1 U9091 ( .A1(n14612), .A2(n14613), .A3(n14614), .A4(n14615), .ZN(
        n14611) );
  NOR2_X1 U9090 ( .A1(n14611), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N146 ) );
  AOI22_X1 U9209 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[31][7] ), .A2(n17154), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[30][7] ), .B2(n17683), .ZN(n14728) );
  AOI22_X1 U9208 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[29][7] ), .A2(n17684), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[28][7] ), .B2(n17685), .ZN(n14729) );
  AOI222_X1 U9207 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[4][7] ), .A2(n17686), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[25][7] ), .B2(n17153), .C1(
        \pipeline/RegFile_DEC_WB/RegBank[24][7] ), .C2(n17687), .ZN(n14730) );
  AOI22_X1 U9206 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[27][7] ), .A2(n17688), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[26][7] ), .B2(n17689), .ZN(n14724) );
  AOI22_X1 U9205 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[23][7] ), .A2(n17690), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[22][7] ), .B2(n17691), .ZN(n14725) );
  AOI22_X1 U9204 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[21][7] ), .A2(n14235), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[20][7] ), .B2(n17693), .ZN(n14726) );
  AOI22_X1 U9203 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[19][7] ), .A2(n17694), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[18][7] ), .B2(n14234), .ZN(n14727) );
  NAND4_X1 U9202 ( .A1(n14724), .A2(n14725), .A3(n14726), .A4(n14727), .ZN(
        n14713) );
  AOI22_X1 U9201 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[17][7] ), .A2(n17696), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[16][7] ), .B2(n17697), .ZN(n14720) );
  AOI22_X1 U9200 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[12][7] ), .A2(n14225), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[13][7] ), .B2(n17358), .ZN(n14721) );
  AOI22_X1 U9199 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[8][7] ), .A2(n17417), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[15][7] ), .B2(n17152), .ZN(n14722) );
  AOI22_X1 U9198 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[9][7] ), .A2(n17352), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[10][7] ), .B2(n14222), .ZN(n14723) );
  NAND4_X1 U9197 ( .A1(n14720), .A2(n14721), .A3(n14722), .A4(n14723), .ZN(
        n14714) );
  AOI22_X1 U9196 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[11][7] ), .A2(n17151), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[3][7] ), .B2(n17413), .ZN(n14716)
         );
  AOI22_X1 U9195 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[14][7] ), .A2(n17700), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[5][7] ), .B2(n17414), .ZN(n14717)
         );
  AOI22_X1 U9194 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[2][7] ), .A2(n17355), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[7][7] ), .B2(n17415), .ZN(n14718)
         );
  AOI22_X1 U9193 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[6][7] ), .A2(n17356), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[1][7] ), .B2(n17416), .ZN(n14719)
         );
  NAND4_X1 U9192 ( .A1(n14716), .A2(n14717), .A3(n14718), .A4(n14719), .ZN(
        n14715) );
  NOR4_X1 U9191 ( .A1(n14712), .A2(n14713), .A3(n14714), .A4(n14715), .ZN(
        n14711) );
  NOR2_X1 U9190 ( .A1(n14711), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N141 ) );
  AOI22_X1 U9129 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[31][11] ), .A2(n17154), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[30][11] ), .B2(n17683), .ZN(
        n14648) );
  AOI22_X1 U9128 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[29][11] ), .A2(n14247), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[28][11] ), .B2(n17685), .ZN(
        n14649) );
  AOI222_X1 U9127 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[4][11] ), .A2(n17686), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[25][11] ), .B2(n17153), .C1(
        \pipeline/RegFile_DEC_WB/RegBank[24][11] ), .C2(n17687), .ZN(n14650)
         );
  AOI22_X1 U9126 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[27][11] ), .A2(n17688), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[26][11] ), .B2(n17689), .ZN(
        n14644) );
  AOI22_X1 U9125 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[23][11] ), .A2(n14237), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[22][11] ), .B2(n17691), .ZN(
        n14645) );
  AOI22_X1 U9124 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[21][11] ), .A2(n17692), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[20][11] ), .B2(n17693), .ZN(
        n14646) );
  AOI22_X1 U9123 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[19][11] ), .A2(n14233), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[18][11] ), .B2(n17695), .ZN(
        n14647) );
  NAND4_X1 U9122 ( .A1(n14644), .A2(n14645), .A3(n14646), .A4(n14647), .ZN(
        n14633) );
  AOI22_X1 U9121 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[17][11] ), .A2(n17696), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[16][11] ), .B2(n17697), .ZN(
        n14640) );
  AOI22_X1 U9120 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[12][11] ), .A2(n17698), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[13][11] ), .B2(n17358), .ZN(
        n14641) );
  AOI22_X1 U9119 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[8][11] ), .A2(n14223), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[15][11] ), .B2(n17152), .ZN(
        n14642) );
  AOI22_X1 U9118 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[9][11] ), .A2(n17352), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[10][11] ), .B2(n17699), .ZN(
        n14643) );
  NAND4_X1 U9117 ( .A1(n14640), .A2(n14641), .A3(n14642), .A4(n14643), .ZN(
        n14634) );
  AOI22_X1 U9116 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[11][11] ), .A2(n17151), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[3][11] ), .B2(n14216), .ZN(n14636) );
  AOI22_X1 U9115 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[14][11] ), .A2(n17700), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[5][11] ), .B2(n14214), .ZN(n14637) );
  AOI22_X1 U9114 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[2][11] ), .A2(n17355), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[7][11] ), .B2(n14212), .ZN(n14638) );
  AOI22_X1 U9113 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[6][11] ), .A2(n17356), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[1][11] ), .B2(n14210), .ZN(n14639) );
  NAND4_X1 U9112 ( .A1(n14636), .A2(n14637), .A3(n14638), .A4(n14639), .ZN(
        n14635) );
  NOR4_X1 U9111 ( .A1(n14632), .A2(n14633), .A3(n14634), .A4(n14635), .ZN(
        n14631) );
  NOR2_X1 U9110 ( .A1(n14631), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N145 ) );
  AOI22_X1 U8769 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[31][29] ), .A2(n17154), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[30][29] ), .B2(n17683), .ZN(
        n14288) );
  AOI22_X1 U8768 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[29][29] ), .A2(n17684), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[28][29] ), .B2(n17685), .ZN(
        n14289) );
  AOI222_X1 U8767 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[4][29] ), .A2(n17686), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[25][29] ), .B2(n17153), .C1(
        \pipeline/RegFile_DEC_WB/RegBank[24][29] ), .C2(n17687), .ZN(n14290)
         );
  AOI22_X1 U8766 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[27][29] ), .A2(n17688), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[26][29] ), .B2(n17689), .ZN(
        n14284) );
  AOI22_X1 U8765 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[23][29] ), .A2(n14237), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[22][29] ), .B2(n17691), .ZN(
        n14285) );
  AOI22_X1 U8764 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[21][29] ), .A2(n17692), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[20][29] ), .B2(n17693), .ZN(
        n14286) );
  AOI22_X1 U8763 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[19][29] ), .A2(n17694), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[18][29] ), .B2(n17695), .ZN(
        n14287) );
  NAND4_X1 U8762 ( .A1(n14284), .A2(n14285), .A3(n14286), .A4(n14287), .ZN(
        n14273) );
  AOI22_X1 U8761 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[17][29] ), .A2(n17696), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[16][29] ), .B2(n17697), .ZN(
        n14280) );
  AOI22_X1 U8760 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[12][29] ), .A2(n17698), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[13][29] ), .B2(n17358), .ZN(
        n14281) );
  AOI22_X1 U8759 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[8][29] ), .A2(n17417), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[15][29] ), .B2(n17152), .ZN(
        n14282) );
  AOI22_X1 U8758 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[9][29] ), .A2(n17352), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[10][29] ), .B2(n17699), .ZN(
        n14283) );
  NAND4_X1 U8757 ( .A1(n14280), .A2(n14281), .A3(n14282), .A4(n14283), .ZN(
        n14274) );
  AOI22_X1 U8756 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[11][29] ), .A2(n17151), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[3][29] ), .B2(n17413), .ZN(n14276) );
  AOI22_X1 U8755 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[14][29] ), .A2(n17700), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[5][29] ), .B2(n17414), .ZN(n14277) );
  AOI22_X1 U8754 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[2][29] ), .A2(n17355), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[7][29] ), .B2(n17415), .ZN(n14278) );
  AOI22_X1 U8753 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[6][29] ), .A2(n17356), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[1][29] ), .B2(n17416), .ZN(n14279) );
  NAND4_X1 U8752 ( .A1(n14276), .A2(n14277), .A3(n14278), .A4(n14279), .ZN(
        n14275) );
  NOR4_X1 U8751 ( .A1(n14272), .A2(n14273), .A3(n14274), .A4(n14275), .ZN(
        n14271) );
  NOR2_X1 U8750 ( .A1(n14271), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N163 ) );
  AOI22_X1 U8749 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[31][30] ), .A2(n17154), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[30][30] ), .B2(n17683), .ZN(
        n14268) );
  AOI22_X1 U8748 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[29][30] ), .A2(n14247), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[28][30] ), .B2(n17685), .ZN(
        n14269) );
  AOI222_X1 U8747 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[4][30] ), .A2(n17686), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[25][30] ), .B2(n17153), .C1(
        \pipeline/RegFile_DEC_WB/RegBank[24][30] ), .C2(n17687), .ZN(n14270)
         );
  AOI22_X1 U8746 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[27][30] ), .A2(n17688), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[26][30] ), .B2(n17689), .ZN(
        n14264) );
  AOI22_X1 U8745 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[23][30] ), .A2(n17690), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[22][30] ), .B2(n17691), .ZN(
        n14265) );
  AOI22_X1 U8744 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[21][30] ), .A2(n17692), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[20][30] ), .B2(n17693), .ZN(
        n14266) );
  AOI22_X1 U8743 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[19][30] ), .A2(n17694), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[18][30] ), .B2(n17695), .ZN(
        n14267) );
  NAND4_X1 U8742 ( .A1(n14264), .A2(n14265), .A3(n14266), .A4(n14267), .ZN(
        n14253) );
  AOI22_X1 U8741 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[17][30] ), .A2(n17696), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[16][30] ), .B2(n17697), .ZN(
        n14260) );
  AOI22_X1 U8740 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[12][30] ), .A2(n17698), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[13][30] ), .B2(n17358), .ZN(
        n14261) );
  AOI22_X1 U8739 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[8][30] ), .A2(n17417), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[15][30] ), .B2(n17152), .ZN(
        n14262) );
  AOI22_X1 U8738 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[9][30] ), .A2(n17352), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[10][30] ), .B2(n17699), .ZN(
        n14263) );
  NAND4_X1 U8737 ( .A1(n14260), .A2(n14261), .A3(n14262), .A4(n14263), .ZN(
        n14254) );
  AOI22_X1 U8736 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[11][30] ), .A2(n17151), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[3][30] ), .B2(n17413), .ZN(n14256) );
  AOI22_X1 U8735 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[14][30] ), .A2(n17700), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[5][30] ), .B2(n17414), .ZN(n14257) );
  AOI22_X1 U8734 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[2][30] ), .A2(n17355), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[7][30] ), .B2(n17415), .ZN(n14258) );
  AOI22_X1 U8733 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[6][30] ), .A2(n17356), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[1][30] ), .B2(n17416), .ZN(n14259) );
  NAND4_X1 U8732 ( .A1(n14256), .A2(n14257), .A3(n14258), .A4(n14259), .ZN(
        n14255) );
  NOR4_X1 U8731 ( .A1(n14252), .A2(n14253), .A3(n14254), .A4(n14255), .ZN(
        n14251) );
  NOR2_X1 U8730 ( .A1(n14251), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N164 ) );
  AOI22_X1 U8849 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[31][25] ), .A2(n17154), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[30][25] ), .B2(n17683), .ZN(
        n14368) );
  AOI22_X1 U8848 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[29][25] ), .A2(n17684), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[28][25] ), .B2(n17685), .ZN(
        n14369) );
  AOI222_X1 U8847 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[4][25] ), .A2(n17686), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[25][25] ), .B2(n17153), .C1(
        \pipeline/RegFile_DEC_WB/RegBank[24][25] ), .C2(n17687), .ZN(n14370)
         );
  AOI22_X1 U8846 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[27][25] ), .A2(n17688), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[26][25] ), .B2(n17689), .ZN(
        n14364) );
  AOI22_X1 U8845 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[23][25] ), .A2(n17690), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[22][25] ), .B2(n17691), .ZN(
        n14365) );
  AOI22_X1 U8844 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[21][25] ), .A2(n17692), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[20][25] ), .B2(n17693), .ZN(
        n14366) );
  AOI22_X1 U8843 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[19][25] ), .A2(n17694), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[18][25] ), .B2(n17695), .ZN(
        n14367) );
  NAND4_X1 U8842 ( .A1(n14364), .A2(n14365), .A3(n14366), .A4(n14367), .ZN(
        n14353) );
  AOI22_X1 U8841 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[17][25] ), .A2(n17696), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[16][25] ), .B2(n17697), .ZN(
        n14360) );
  AOI22_X1 U8840 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[12][25] ), .A2(n17698), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[13][25] ), .B2(n17357), .ZN(
        n14361) );
  AOI22_X1 U8839 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[8][25] ), .A2(n17417), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[15][25] ), .B2(n17152), .ZN(
        n14362) );
  AOI22_X1 U8838 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[9][25] ), .A2(n17351), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[10][25] ), .B2(n17699), .ZN(
        n14363) );
  NAND4_X1 U8837 ( .A1(n14360), .A2(n14361), .A3(n14362), .A4(n14363), .ZN(
        n14354) );
  AOI22_X1 U8836 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[11][25] ), .A2(n17151), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[3][25] ), .B2(n17413), .ZN(n14356) );
  AOI22_X1 U8835 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[14][25] ), .A2(n17700), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[5][25] ), .B2(n17414), .ZN(n14357) );
  AOI22_X1 U8834 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[2][25] ), .A2(n17353), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[7][25] ), .B2(n17415), .ZN(n14358) );
  AOI22_X1 U8833 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[6][25] ), .A2(n17354), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[1][25] ), .B2(n17416), .ZN(n14359) );
  NAND4_X1 U8832 ( .A1(n14356), .A2(n14357), .A3(n14358), .A4(n14359), .ZN(
        n14355) );
  NOR4_X1 U8831 ( .A1(n14352), .A2(n14353), .A3(n14354), .A4(n14355), .ZN(
        n14351) );
  NOR2_X1 U8830 ( .A1(n14351), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N159 ) );
  AOI22_X1 U9289 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[31][3] ), .A2(n17154), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[30][3] ), .B2(n17683), .ZN(n14808) );
  AOI22_X1 U9288 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[29][3] ), .A2(n14247), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[28][3] ), .B2(n17685), .ZN(n14809) );
  AOI222_X1 U9287 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[4][3] ), .A2(n17686), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[25][3] ), .B2(n17153), .C1(
        \pipeline/RegFile_DEC_WB/RegBank[24][3] ), .C2(n17687), .ZN(n14810) );
  AOI22_X1 U9286 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[27][3] ), .A2(n17688), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[26][3] ), .B2(n17689), .ZN(n14804) );
  AOI22_X1 U9285 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[23][3] ), .A2(n17690), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[22][3] ), .B2(n17691), .ZN(n14805) );
  AOI22_X1 U9284 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[21][3] ), .A2(n17692), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[20][3] ), .B2(n17693), .ZN(n14806) );
  AOI22_X1 U9283 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[19][3] ), .A2(n14233), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[18][3] ), .B2(n17695), .ZN(n14807) );
  NAND4_X1 U9282 ( .A1(n14804), .A2(n14805), .A3(n14806), .A4(n14807), .ZN(
        n14793) );
  AOI22_X1 U9281 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[17][3] ), .A2(n17696), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[16][3] ), .B2(n17697), .ZN(n14800) );
  AOI22_X1 U9280 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[12][3] ), .A2(n17698), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[13][3] ), .B2(n17357), .ZN(n14801) );
  AOI22_X1 U9279 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[8][3] ), .A2(n17417), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[15][3] ), .B2(n17152), .ZN(n14802) );
  AOI22_X1 U9278 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[9][3] ), .A2(n17351), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[10][3] ), .B2(n17699), .ZN(n14803) );
  NAND4_X1 U9277 ( .A1(n14800), .A2(n14801), .A3(n14802), .A4(n14803), .ZN(
        n14794) );
  AOI22_X1 U9276 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[11][3] ), .A2(n17151), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[3][3] ), .B2(n17413), .ZN(n14796)
         );
  AOI22_X1 U9275 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[14][3] ), .A2(n17700), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[5][3] ), .B2(n17414), .ZN(n14797)
         );
  AOI22_X1 U9274 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[2][3] ), .A2(n17353), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[7][3] ), .B2(n17415), .ZN(n14798)
         );
  AOI22_X1 U9273 ( .A1(\pipeline/RegFile_DEC_WB/RegBank[6][3] ), .A2(n17354), 
        .B1(\pipeline/RegFile_DEC_WB/RegBank[1][3] ), .B2(n17416), .ZN(n14799)
         );
  NAND4_X1 U9272 ( .A1(n14796), .A2(n14797), .A3(n14798), .A4(n14799), .ZN(
        n14795) );
  NOR4_X1 U9271 ( .A1(n14792), .A2(n14793), .A3(n14794), .A4(n14795), .ZN(
        n14791) );
  NOR2_X1 U9270 ( .A1(n14791), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N137 ) );
  OAI22_X1 U9420 ( .A1(n14913), .A2(n17075), .B1(n17109), .B2(n17461), .ZN(
        \pipeline/IDEX_Stage/N118 ) );
  OAI22_X1 U9402 ( .A1(n14895), .A2(n17075), .B1(n17682), .B2(n17451), .ZN(
        \pipeline/IDEX_Stage/N127 ) );
  OAI22_X1 U9452 ( .A1(n14945), .A2(n17075), .B1(n17109), .B2(n17450), .ZN(
        \pipeline/IDEX_Stage/N102 ) );
  OAI22_X1 U9442 ( .A1(n14935), .A2(n17075), .B1(n17109), .B2(n17454), .ZN(
        \pipeline/IDEX_Stage/N107 ) );
  OAI22_X1 U9414 ( .A1(n14907), .A2(n17075), .B1(n17109), .B2(n17438), .ZN(
        \pipeline/IDEX_Stage/N121 ) );
  OAI22_X1 U9390 ( .A1(n14883), .A2(n17075), .B1(n17109), .B2(n17527), .ZN(
        \pipeline/IDEX_Stage/N133 ) );
  NOR2_X1 U8698 ( .A1(n17350), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N171 ) );
  NOR2_X1 U8668 ( .A1(n17349), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N206 ) );
  NOR2_X1 U8686 ( .A1(n17433), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N177 ) );
  NOR2_X1 U8696 ( .A1(n17361), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N172 ) );
  NOR2_X1 U8702 ( .A1(n17410), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N169 ) );
  NOR2_X1 U8706 ( .A1(n17406), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N167 ) );
  NOR2_X1 U8684 ( .A1(n17444), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N178 ) );
  NOR2_X1 U8674 ( .A1(n17383), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N200 ) );
  NOR2_X1 U8694 ( .A1(n17437), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N173 ) );
  NOR2_X1 U8669 ( .A1(n17408), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N205 ) );
  NOR2_X1 U8672 ( .A1(n17328), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N202 ) );
  NOR2_X1 U8673 ( .A1(n17384), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N201 ) );
  NOR2_X1 U8671 ( .A1(n17316), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N203 ) );
  OAI22_X1 U9394 ( .A1(n14887), .A2(n17075), .B1(n17109), .B2(n17452), .ZN(
        \pipeline/IDEX_Stage/N131 ) );
  OAI22_X1 U9422 ( .A1(n14915), .A2(n17075), .B1(n17109), .B2(n17453), .ZN(
        \pipeline/IDEX_Stage/N117 ) );
  OAI22_X1 U9424 ( .A1(n14917), .A2(n17075), .B1(n17682), .B2(n17460), .ZN(
        \pipeline/IDEX_Stage/N116 ) );
  NOR2_X1 U8690 ( .A1(n17432), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N175 ) );
  NOR2_X1 U8675 ( .A1(n17317), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N199 ) );
  NOR2_X1 U8708 ( .A1(n17076), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N166 ) );
  NOR2_X1 U8682 ( .A1(n17434), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N179 ) );
  NOR2_X1 U8692 ( .A1(n17428), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N174 ) );
  NOR2_X1 U8680 ( .A1(n17445), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N180 ) );
  NOR2_X1 U8700 ( .A1(n17412), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N170 ) );
  NOR2_X1 U8670 ( .A1(n17329), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N204 ) );
  NOR2_X1 U8667 ( .A1(n17407), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N207 ) );
  NOR2_X1 U8676 ( .A1(n17315), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N198 ) );
  NOR2_X1 U8688 ( .A1(n17440), .A2(n17075), .ZN(\pipeline/IDEX_Stage/N176 ) );
  AOI22_X1 U8594 ( .A1(\pipeline/Alu_Out_Addr_to_mem[1] ), .A2(n17370), .B1(
        n14135), .B2(data_from_dram[1]), .ZN(n14165) );
  AOI22_X1 U8596 ( .A1(\pipeline/Alu_Out_Addr_to_mem[0] ), .A2(n17370), .B1(
        n14135), .B2(data_from_dram[0]), .ZN(n14166) );
  AOI22_X1 U8566 ( .A1(\pipeline/Alu_Out_Addr_to_mem[15] ), .A2(n14134), .B1(
        n14135), .B2(data_from_dram[15]), .ZN(n14151) );
  AOI22_X1 U8570 ( .A1(\pipeline/Alu_Out_Addr_to_mem[13] ), .A2(n14134), .B1(
        n14135), .B2(data_from_dram[13]), .ZN(n14153) );
  AOI22_X1 U8548 ( .A1(\pipeline/Alu_Out_Addr_to_mem[24] ), .A2(n17370), .B1(
        n14135), .B2(data_from_dram[24]), .ZN(n14142) );
  AOI22_X1 U8584 ( .A1(\pipeline/Alu_Out_Addr_to_mem[6] ), .A2(n17370), .B1(
        n14135), .B2(data_from_dram[6]), .ZN(n14160) );
  AOI22_X1 U8540 ( .A1(\pipeline/Alu_Out_Addr_to_mem[28] ), .A2(n17370), .B1(
        n14135), .B2(data_from_dram[28]), .ZN(n14138) );
  AOI22_X1 U8572 ( .A1(\pipeline/Alu_Out_Addr_to_mem[12] ), .A2(n14134), .B1(
        n14135), .B2(data_from_dram[12]), .ZN(n14154) );
  AOI22_X1 U8534 ( .A1(\pipeline/Alu_Out_Addr_to_mem[31] ), .A2(n14134), .B1(
        n14135), .B2(data_from_dram[31]), .ZN(n14133) );
  AOI22_X1 U8546 ( .A1(\pipeline/Alu_Out_Addr_to_mem[25] ), .A2(n17370), .B1(
        n14135), .B2(data_from_dram[25]), .ZN(n14141) );
  AOI22_X1 U8550 ( .A1(\pipeline/Alu_Out_Addr_to_mem[23] ), .A2(n17370), .B1(
        n14135), .B2(data_from_dram[23]), .ZN(n14143) );
  AOI22_X1 U8588 ( .A1(\pipeline/Alu_Out_Addr_to_mem[4] ), .A2(n17370), .B1(
        n14135), .B2(data_from_dram[4]), .ZN(n14162) );
  AOI22_X1 U8590 ( .A1(\pipeline/Alu_Out_Addr_to_mem[3] ), .A2(n17370), .B1(
        n14135), .B2(data_from_dram[3]), .ZN(n14163) );
  AOI22_X1 U8580 ( .A1(\pipeline/Alu_Out_Addr_to_mem[8] ), .A2(n17370), .B1(
        n14135), .B2(data_from_dram[8]), .ZN(n14158) );
  AOI22_X1 U8582 ( .A1(\pipeline/Alu_Out_Addr_to_mem[7] ), .A2(n17370), .B1(
        n14135), .B2(data_from_dram[7]), .ZN(n14159) );
  AOI22_X1 U8552 ( .A1(\pipeline/Alu_Out_Addr_to_mem[22] ), .A2(n17370), .B1(
        n14135), .B2(data_from_dram[22]), .ZN(n14144) );
  AOI22_X1 U8592 ( .A1(\pipeline/Alu_Out_Addr_to_mem[2] ), .A2(n17370), .B1(
        n14135), .B2(data_from_dram[2]), .ZN(n14164) );
  AOI22_X1 U8578 ( .A1(\pipeline/Alu_Out_Addr_to_mem[9] ), .A2(n14134), .B1(
        n14135), .B2(data_from_dram[9]), .ZN(n14157) );
  AOI22_X1 U8554 ( .A1(\pipeline/Alu_Out_Addr_to_mem[21] ), .A2(n14134), .B1(
        n14135), .B2(data_from_dram[21]), .ZN(n14145) );
  AOI22_X1 U8574 ( .A1(\pipeline/Alu_Out_Addr_to_mem[11] ), .A2(n14134), .B1(
        n14135), .B2(data_from_dram[11]), .ZN(n14155) );
  AOI22_X1 U8560 ( .A1(\pipeline/Alu_Out_Addr_to_mem[18] ), .A2(n14134), .B1(
        n14135), .B2(data_from_dram[18]), .ZN(n14148) );
  AOI22_X1 U8556 ( .A1(\pipeline/Alu_Out_Addr_to_mem[20] ), .A2(n14134), .B1(
        n14135), .B2(data_from_dram[20]), .ZN(n14146) );
  AOI22_X1 U8536 ( .A1(\pipeline/Alu_Out_Addr_to_mem[30] ), .A2(n17370), .B1(
        n14135), .B2(data_from_dram[30]), .ZN(n14136) );
  AOI22_X1 U8538 ( .A1(\pipeline/Alu_Out_Addr_to_mem[29] ), .A2(n17370), .B1(
        n14135), .B2(data_from_dram[29]), .ZN(n14137) );
  AOI22_X1 U8542 ( .A1(\pipeline/Alu_Out_Addr_to_mem[27] ), .A2(n17370), .B1(
        n14135), .B2(data_from_dram[27]), .ZN(n14139) );
  AOI22_X1 U8558 ( .A1(\pipeline/Alu_Out_Addr_to_mem[19] ), .A2(n14134), .B1(
        n14135), .B2(data_from_dram[19]), .ZN(n14147) );
  AOI22_X1 U8544 ( .A1(\pipeline/Alu_Out_Addr_to_mem[26] ), .A2(n17370), .B1(
        n14135), .B2(data_from_dram[26]), .ZN(n14140) );
  AOI22_X1 U8568 ( .A1(\pipeline/Alu_Out_Addr_to_mem[14] ), .A2(n14134), .B1(
        n14135), .B2(data_from_dram[14]), .ZN(n14152) );
  AOI22_X1 U8586 ( .A1(\pipeline/Alu_Out_Addr_to_mem[5] ), .A2(n17370), .B1(
        n14135), .B2(data_from_dram[5]), .ZN(n14161) );
  AOI22_X1 U8562 ( .A1(\pipeline/Alu_Out_Addr_to_mem[17] ), .A2(n14134), .B1(
        n14135), .B2(data_from_dram[17]), .ZN(n14149) );
  AOI22_X1 U8564 ( .A1(\pipeline/Alu_Out_Addr_to_mem[16] ), .A2(n14134), .B1(
        n14135), .B2(data_from_dram[16]), .ZN(n14150) );
  AOI22_X1 U8576 ( .A1(\pipeline/Alu_Out_Addr_to_mem[10] ), .A2(n14134), .B1(
        n14135), .B2(data_from_dram[10]), .ZN(n14156) );
  NAND2_X1 U8608 ( .A1(n17703), .A2(n14007), .ZN(n13988) );
  NOR2_X1 U8607 ( .A1(n14168), .A2(n13988), .ZN(\pipeline/IDEX_Stage/N92 ) );
  NOR2_X1 U8611 ( .A1(n17382), .A2(n14169), .ZN(n14123) );
  NOR2_X1 U8609 ( .A1(n14168), .A2(n13981), .ZN(\pipeline/IDEX_Stage/N91 ) );
  AOI21_X1 U8663 ( .B1(n14025), .B2(n17349), .A(n14168), .ZN(
        \pipeline/IDEX_Stage/N211 ) );
  AOI21_X1 U8704 ( .B1(n14025), .B2(n17404), .A(n14168), .ZN(
        \pipeline/IDEX_Stage/N168 ) );
  AOI21_X1 U8664 ( .B1(n14025), .B2(n17408), .A(n14168), .ZN(
        \pipeline/IDEX_Stage/N210 ) );
  AOI21_X1 U8659 ( .B1(n14025), .B2(n17434), .A(n14168), .ZN(
        \pipeline/IDEX_Stage/N215 ) );
  AOI21_X1 U8657 ( .B1(n14025), .B2(n17431), .A(n14168), .ZN(
        \pipeline/IDEX_Stage/N217 ) );
  AOI21_X1 U8658 ( .B1(n14025), .B2(n17445), .A(n14168), .ZN(
        \pipeline/IDEX_Stage/N216 ) );
  AOI21_X1 U8662 ( .B1(n14025), .B2(n17407), .A(n14168), .ZN(
        \pipeline/IDEX_Stage/N212 ) );
  AOI21_X1 U8666 ( .B1(n14025), .B2(n17316), .A(n14168), .ZN(
        \pipeline/IDEX_Stage/N208 ) );
  AOI21_X1 U8665 ( .B1(n14025), .B2(n17329), .A(n14168), .ZN(
        \pipeline/IDEX_Stage/N209 ) );
  AOI21_X1 U8660 ( .B1(n14025), .B2(n17444), .A(n14168), .ZN(
        \pipeline/IDEX_Stage/N214 ) );
  AOI21_X1 U8661 ( .B1(n14025), .B2(n17433), .A(n14168), .ZN(
        \pipeline/IDEX_Stage/N213 ) );
  NOR3_X1 U9474 ( .A1(n14982), .A2(n17447), .A3(n14129), .ZN(
        \pipeline/EXMEM_stage/N76 ) );
  NOR2_X1 U8528 ( .A1(n17393), .A2(n14129), .ZN(\pipeline/MEMWB_Stage/N47 ) );
  NOR2_X1 U8531 ( .A1(n17645), .A2(n14129), .ZN(\pipeline/MEMWB_Stage/N44 ) );
  NOR2_X1 U8530 ( .A1(n17646), .A2(n14129), .ZN(\pipeline/MEMWB_Stage/N45 ) );
  NOR2_X1 U9476 ( .A1(n13281), .A2(n14101), .ZN(\pipeline/EXMEM_stage/N75 ) );
  AOI22_X1 U9483 ( .A1(\pipeline/EXE_controls_in_EXEcute [7]), .A2(n13931), 
        .B1(n13926), .B2(n17430), .ZN(n14117) );
  NOR2_X1 U9482 ( .A1(n13281), .A2(n14117), .ZN(\pipeline/EXMEM_stage/N72 ) );
  AOI22_X1 U9485 ( .A1(\pipeline/EXE_controls_in_EXEcute [7]), .A2(n13930), 
        .B1(n13925), .B2(n17430), .ZN(n14116) );
  NOR2_X1 U9484 ( .A1(n13281), .A2(n14116), .ZN(\pipeline/EXMEM_stage/N71 ) );
  OAI21_X1 U10044 ( .B1(n15646), .B2(n17371), .A(n17703), .ZN(n3925) );
  OAI21_X1 U10042 ( .B1(n15646), .B2(n17372), .A(n17703), .ZN(n3926) );
  OAI21_X1 U10022 ( .B1(n15646), .B2(n17478), .A(n17702), .ZN(n3936) );
  OAI21_X1 U10038 ( .B1(n15646), .B2(n17472), .A(n17702), .ZN(n3928) );
  OAI21_X1 U10016 ( .B1(n15646), .B2(n17481), .A(n17702), .ZN(n3939) );
  OAI21_X1 U10018 ( .B1(n15646), .B2(n17480), .A(n17702), .ZN(n3938) );
  OAI21_X1 U10020 ( .B1(n15646), .B2(n17479), .A(n17702), .ZN(n3937) );
  OAI21_X1 U10026 ( .B1(n15646), .B2(n17477), .A(n17702), .ZN(n3934) );
  OAI21_X1 U10028 ( .B1(n15646), .B2(n17476), .A(n17702), .ZN(n3933) );
  OAI21_X1 U10024 ( .B1(n15646), .B2(n17375), .A(n17701), .ZN(n3935) );
  OAI21_X1 U10004 ( .B1(n15646), .B2(n17378), .A(n17701), .ZN(n3945) );
  OAI21_X1 U10002 ( .B1(n15646), .B2(n17485), .A(n17701), .ZN(n3946) );
  OAI21_X1 U10000 ( .B1(n15646), .B2(n17486), .A(n17701), .ZN(n3947) );
  OAI21_X1 U9998 ( .B1(n15646), .B2(n17487), .A(n17701), .ZN(n3948) );
  OAI21_X1 U9996 ( .B1(n15646), .B2(n17488), .A(n17701), .ZN(n3949) );
  OAI21_X1 U9994 ( .B1(n15646), .B2(n17489), .A(n17701), .ZN(n3950) );
  OAI21_X1 U9992 ( .B1(n15646), .B2(n17490), .A(n17701), .ZN(n3951) );
  OAI21_X1 U9990 ( .B1(n15646), .B2(n17491), .A(n17701), .ZN(n3952) );
  OAI21_X1 U10014 ( .B1(n15646), .B2(n17376), .A(n17702), .ZN(n3940) );
  OAI21_X1 U10012 ( .B1(n15646), .B2(n17377), .A(n17701), .ZN(n3941) );
  OAI21_X1 U10010 ( .B1(n15646), .B2(n17482), .A(n17701), .ZN(n3942) );
  OAI21_X1 U10008 ( .B1(n15646), .B2(n17483), .A(n17701), .ZN(n3943) );
  OAI21_X1 U10006 ( .B1(n15646), .B2(n17484), .A(n17701), .ZN(n3944) );
  OAI21_X1 U10030 ( .B1(n15646), .B2(n17475), .A(n17702), .ZN(n3932) );
  OAI21_X1 U10032 ( .B1(n15646), .B2(n17474), .A(n17702), .ZN(n3931) );
  OAI21_X1 U10034 ( .B1(n15646), .B2(n17473), .A(n17702), .ZN(n3930) );
  OAI21_X1 U10036 ( .B1(n15646), .B2(n17374), .A(n17702), .ZN(n3929) );
  OAI21_X1 U10040 ( .B1(n15646), .B2(n17373), .A(n17702), .ZN(n3927) );
  AOI22_X1 U9481 ( .A1(\pipeline/EXE_controls_in_EXEcute [7]), .A2(n13932), 
        .B1(n13927), .B2(n17430), .ZN(n14113) );
  NOR2_X1 U9480 ( .A1(n13281), .A2(n14113), .ZN(\pipeline/EXMEM_stage/N73 ) );
  AOI22_X1 U9479 ( .A1(\pipeline/EXE_controls_in_EXEcute [7]), .A2(n13933), 
        .B1(n13928), .B2(n17430), .ZN(n14100) );
  NOR2_X1 U9478 ( .A1(n13281), .A2(n14100), .ZN(\pipeline/EXMEM_stage/N74 ) );
  OAI21_X1 U9984 ( .B1(n15646), .B2(n17494), .A(n17701), .ZN(n3955) );
  OAI21_X1 U9982 ( .B1(n15646), .B2(n17379), .A(n17702), .ZN(n3956) );
  OAI21_X1 U9986 ( .B1(n15646), .B2(n17493), .A(n17702), .ZN(n3954) );
  OAI21_X1 U9988 ( .B1(n15646), .B2(n17492), .A(n17705), .ZN(n3953) );
  NOR2_X1 U9563 ( .A1(n13281), .A2(n17447), .ZN(\pipeline/EXMEM_stage/N5 ) );
  NOR2_X1 U9585 ( .A1(n13281), .A2(n17449), .ZN(\pipeline/EXMEM_stage/N4 ) );
  OAI21_X1 U11058 ( .B1(n15001), .B2(n16598), .A(
        \pipeline/EXE_controls_in_EXEcute [5]), .ZN(n16599) );
  AOI211_X1 U11057 ( .C1(n15001), .C2(n16598), .A(
        \pipeline/EXE_controls_in_EXEcute [6]), .B(n16599), .ZN(exception) );
  NOR2_X1 U11949 ( .A1(n17000), .A2(n16597), .ZN(\DataMem/N1671 ) );
  NOR2_X1 U11894 ( .A1(n17000), .A2(n16596), .ZN(\DataMem/N1735 ) );
  NOR2_X1 U11859 ( .A1(n17000), .A2(n16595), .ZN(\DataMem/N1799 ) );
  AOI22_X1 U11599 ( .A1(n16823), .A2(\DataMem/Mem[7][11] ), .B1(n16824), .B2(
        \DataMem/Mem[6][11] ), .ZN(n16921) );
  NAND2_X1 U11769 ( .A1(addr_to_dataRam[4]), .A2(addr_to_dataRam[2]), .ZN(
        n17014) );
  AOI22_X1 U11598 ( .A1(n16821), .A2(\DataMem/Mem[5][11] ), .B1(n16822), .B2(
        \DataMem/Mem[4][11] ), .ZN(n16922) );
  NAND2_X1 U11838 ( .A1(addr_to_dataRam[2]), .A2(addr_to_dataRam[3]), .ZN(
        n17016) );
  NOR3_X1 U11872 ( .A1(addr_to_dataRam[4]), .A2(addr_to_dataRam[2]), .A3(
        n17015), .ZN(n16820) );
  AOI22_X1 U11597 ( .A1(n17122), .A2(\DataMem/Mem[3][11] ), .B1(n17653), .B2(
        \DataMem/Mem[2][11] ), .ZN(n16923) );
  AOI22_X1 U11596 ( .A1(n17124), .A2(\DataMem/Mem[1][11] ), .B1(n17125), .B2(
        \DataMem/Mem[0][11] ), .ZN(n16924) );
  NOR2_X1 U11594 ( .A1(n17155), .A2(n16920), .ZN(\DataMem/N2194 ) );
  NOR2_X1 U11687 ( .A1(n17001), .A2(n16590), .ZN(\DataMem/N2117 ) );
  NOR2_X1 U11721 ( .A1(n17001), .A2(n16591), .ZN(\DataMem/N2053 ) );
  NOR2_X1 U11756 ( .A1(n17001), .A2(n16592), .ZN(\DataMem/N1989 ) );
  NOR2_X1 U11791 ( .A1(n17001), .A2(n16593), .ZN(\DataMem/N1925 ) );
  NOR2_X1 U11825 ( .A1(n17001), .A2(n16594), .ZN(\DataMem/N1861 ) );
  NOR2_X1 U11860 ( .A1(n17001), .A2(n16595), .ZN(\DataMem/N1797 ) );
  NOR2_X1 U11895 ( .A1(n17001), .A2(n16596), .ZN(\DataMem/N1733 ) );
  NOR2_X1 U11947 ( .A1(n16999), .A2(n17650), .ZN(\DataMem/N1673 ) );
  AOI22_X1 U11593 ( .A1(n16823), .A2(\DataMem/Mem[7][12] ), .B1(n16824), .B2(
        \DataMem/Mem[6][12] ), .ZN(n16916) );
  AOI22_X1 U11592 ( .A1(n16821), .A2(\DataMem/Mem[5][12] ), .B1(n16822), .B2(
        \DataMem/Mem[4][12] ), .ZN(n16917) );
  AOI22_X1 U11591 ( .A1(n17122), .A2(\DataMem/Mem[3][12] ), .B1(n17653), .B2(
        \DataMem/Mem[2][12] ), .ZN(n16918) );
  AOI22_X1 U11590 ( .A1(n17124), .A2(\DataMem/Mem[1][12] ), .B1(n17125), .B2(
        \DataMem/Mem[0][12] ), .ZN(n16919) );
  NOR2_X1 U11588 ( .A1(n17155), .A2(n16915), .ZN(\DataMem/N2197 ) );
  NOR2_X1 U11695 ( .A1(n17009), .A2(n17661), .ZN(\DataMem/N2101 ) );
  NOR2_X1 U11729 ( .A1(n17009), .A2(n17658), .ZN(\DataMem/N2037 ) );
  NOR2_X1 U11764 ( .A1(n17009), .A2(n17657), .ZN(\DataMem/N1973 ) );
  NOR2_X1 U11799 ( .A1(n17009), .A2(n17656), .ZN(\DataMem/N1909 ) );
  NOR2_X1 U11833 ( .A1(n17009), .A2(n17655), .ZN(\DataMem/N1845 ) );
  NOR2_X1 U11868 ( .A1(n17009), .A2(n17654), .ZN(\DataMem/N1781 ) );
  NOR2_X1 U11903 ( .A1(n17009), .A2(n17651), .ZN(\DataMem/N1717 ) );
  NOR2_X1 U11967 ( .A1(n17009), .A2(n17650), .ZN(\DataMem/N1653 ) );
  AOI22_X1 U11940 ( .A1(\pipeline/Forward_sw1_mux ), .A2(
        \pipeline/data_to_RF_from_WB[16] ), .B1(n13803), .B2(n17380), .ZN(
        n16995) );
  NOR2_X1 U11854 ( .A1(n16995), .A2(n17654), .ZN(\DataMem/N1809 ) );
  AOI22_X1 U11653 ( .A1(n17659), .A2(\DataMem/Mem[7][2] ), .B1(n17530), .B2(
        \DataMem/Mem[6][2] ), .ZN(n16966) );
  AOI22_X1 U11652 ( .A1(n17531), .A2(\DataMem/Mem[5][2] ), .B1(n16822), .B2(
        \DataMem/Mem[4][2] ), .ZN(n16967) );
  AOI22_X1 U11651 ( .A1(n17122), .A2(\DataMem/Mem[3][2] ), .B1(n17653), .B2(
        \DataMem/Mem[2][2] ), .ZN(n16968) );
  AOI22_X1 U11650 ( .A1(n17124), .A2(\DataMem/Mem[1][2] ), .B1(n17125), .B2(
        \DataMem/Mem[0][2] ), .ZN(n16969) );
  NOR2_X1 U11648 ( .A1(n17155), .A2(n16965), .ZN(\DataMem/N2167 ) );
  NOR2_X1 U11694 ( .A1(n17008), .A2(n17661), .ZN(\DataMem/N2103 ) );
  NOR2_X1 U11728 ( .A1(n17008), .A2(n17658), .ZN(\DataMem/N2039 ) );
  NOR2_X1 U11763 ( .A1(n17008), .A2(n17657), .ZN(\DataMem/N1975 ) );
  NOR2_X1 U11798 ( .A1(n17008), .A2(n17656), .ZN(\DataMem/N1911 ) );
  NOR2_X1 U11832 ( .A1(n17008), .A2(n17655), .ZN(\DataMem/N1847 ) );
  NOR2_X1 U11867 ( .A1(n17008), .A2(n17654), .ZN(\DataMem/N1783 ) );
  NOR2_X1 U11902 ( .A1(n17008), .A2(n17651), .ZN(\DataMem/N1719 ) );
  NOR2_X1 U11965 ( .A1(n17008), .A2(n17650), .ZN(\DataMem/N1655 ) );
  AOI22_X1 U11647 ( .A1(n17660), .A2(\DataMem/Mem[7][3] ), .B1(n17530), .B2(
        \DataMem/Mem[6][3] ), .ZN(n16961) );
  AOI22_X1 U11646 ( .A1(n17531), .A2(\DataMem/Mem[5][3] ), .B1(n16822), .B2(
        \DataMem/Mem[4][3] ), .ZN(n16962) );
  AOI22_X1 U11645 ( .A1(n17122), .A2(\DataMem/Mem[3][3] ), .B1(n17653), .B2(
        \DataMem/Mem[2][3] ), .ZN(n16963) );
  AOI22_X1 U11644 ( .A1(n17124), .A2(\DataMem/Mem[1][3] ), .B1(n17125), .B2(
        \DataMem/Mem[0][3] ), .ZN(n16964) );
  NOR2_X1 U11642 ( .A1(n17155), .A2(n16960), .ZN(\DataMem/N2170 ) );
  NOR2_X1 U11681 ( .A1(n16995), .A2(n17661), .ZN(\DataMem/N2129 ) );
  NOR2_X1 U11715 ( .A1(n16995), .A2(n17658), .ZN(\DataMem/N2065 ) );
  NOR2_X1 U11750 ( .A1(n16995), .A2(n17657), .ZN(\DataMem/N2001 ) );
  NOR2_X1 U11785 ( .A1(n16995), .A2(n17656), .ZN(\DataMem/N1937 ) );
  NOR2_X1 U11819 ( .A1(n16995), .A2(n17655), .ZN(\DataMem/N1873 ) );
  NOR2_X1 U11685 ( .A1(n16999), .A2(n17661), .ZN(\DataMem/N2121 ) );
  NOR2_X1 U11719 ( .A1(n16999), .A2(n17658), .ZN(\DataMem/N2057 ) );
  NOR2_X1 U11754 ( .A1(n16999), .A2(n17657), .ZN(\DataMem/N1993 ) );
  NOR2_X1 U11789 ( .A1(n16999), .A2(n17656), .ZN(\DataMem/N1929 ) );
  NOR2_X1 U11823 ( .A1(n16999), .A2(n17655), .ZN(\DataMem/N1865 ) );
  NOR2_X1 U11858 ( .A1(n16999), .A2(n17654), .ZN(\DataMem/N1801 ) );
  NOR2_X1 U11893 ( .A1(n16999), .A2(n17651), .ZN(\DataMem/N1737 ) );
  NOR2_X1 U11696 ( .A1(n17010), .A2(n17661), .ZN(\DataMem/N2099 ) );
  NOR2_X1 U11730 ( .A1(n17010), .A2(n17658), .ZN(\DataMem/N2035 ) );
  NOR2_X1 U11765 ( .A1(n17010), .A2(n17657), .ZN(\DataMem/N1971 ) );
  NOR2_X1 U11800 ( .A1(n17010), .A2(n17656), .ZN(\DataMem/N1907 ) );
  NOR2_X1 U11834 ( .A1(n17010), .A2(n17655), .ZN(\DataMem/N1843 ) );
  NOR2_X1 U11869 ( .A1(n17010), .A2(n17654), .ZN(\DataMem/N1779 ) );
  NOR2_X1 U11904 ( .A1(n17010), .A2(n17651), .ZN(\DataMem/N1715 ) );
  NOR2_X1 U11759 ( .A1(n17004), .A2(n17657), .ZN(\DataMem/N1983 ) );
  NOR2_X1 U11693 ( .A1(n17007), .A2(n17661), .ZN(\DataMem/N2105 ) );
  NOR2_X1 U11727 ( .A1(n17007), .A2(n17658), .ZN(\DataMem/N2041 ) );
  NOR2_X1 U11762 ( .A1(n17007), .A2(n17657), .ZN(\DataMem/N1977 ) );
  NOR2_X1 U11797 ( .A1(n17007), .A2(n17656), .ZN(\DataMem/N1913 ) );
  NOR2_X1 U11831 ( .A1(n17007), .A2(n17655), .ZN(\DataMem/N1849 ) );
  NOR2_X1 U11866 ( .A1(n17007), .A2(n17654), .ZN(\DataMem/N1785 ) );
  NOR2_X1 U11901 ( .A1(n17007), .A2(n17651), .ZN(\DataMem/N1721 ) );
  NOR2_X1 U11963 ( .A1(n17007), .A2(n17650), .ZN(\DataMem/N1657 ) );
  AOI22_X1 U11641 ( .A1(n17660), .A2(\DataMem/Mem[7][4] ), .B1(n17530), .B2(
        \DataMem/Mem[6][4] ), .ZN(n16956) );
  AOI22_X1 U11640 ( .A1(n17531), .A2(\DataMem/Mem[5][4] ), .B1(n16822), .B2(
        \DataMem/Mem[4][4] ), .ZN(n16957) );
  AOI22_X1 U11639 ( .A1(n17122), .A2(\DataMem/Mem[3][4] ), .B1(n17652), .B2(
        \DataMem/Mem[2][4] ), .ZN(n16958) );
  AOI22_X1 U11638 ( .A1(n17124), .A2(\DataMem/Mem[1][4] ), .B1(n17125), .B2(
        \DataMem/Mem[0][4] ), .ZN(n16959) );
  NOR2_X1 U11636 ( .A1(n17155), .A2(n16955), .ZN(\DataMem/N2173 ) );
  AOI22_X1 U11605 ( .A1(n16823), .A2(\DataMem/Mem[7][10] ), .B1(n16824), .B2(
        \DataMem/Mem[6][10] ), .ZN(n16926) );
  AOI22_X1 U11604 ( .A1(n16821), .A2(\DataMem/Mem[5][10] ), .B1(n16822), .B2(
        \DataMem/Mem[4][10] ), .ZN(n16927) );
  AOI22_X1 U11603 ( .A1(n17122), .A2(\DataMem/Mem[3][10] ), .B1(n17653), .B2(
        \DataMem/Mem[2][10] ), .ZN(n16928) );
  AOI22_X1 U11602 ( .A1(n17124), .A2(\DataMem/Mem[1][10] ), .B1(n17125), .B2(
        \DataMem/Mem[0][10] ), .ZN(n16929) );
  NOR2_X1 U11600 ( .A1(n17155), .A2(n16925), .ZN(\DataMem/N2191 ) );
  NOR2_X1 U11951 ( .A1(n17001), .A2(n16597), .ZN(\DataMem/N1669 ) );
  NOR2_X1 U11899 ( .A1(n17005), .A2(n17651), .ZN(\DataMem/N1725 ) );
  NOR2_X1 U11864 ( .A1(n17005), .A2(n17654), .ZN(\DataMem/N1789 ) );
  NOR2_X1 U11829 ( .A1(n17005), .A2(n17655), .ZN(\DataMem/N1853 ) );
  NOR2_X1 U11795 ( .A1(n17005), .A2(n17656), .ZN(\DataMem/N1917 ) );
  NOR2_X1 U11760 ( .A1(n17005), .A2(n17657), .ZN(\DataMem/N1981 ) );
  NOR2_X1 U11725 ( .A1(n17005), .A2(n17658), .ZN(\DataMem/N2045 ) );
  NOR2_X1 U11691 ( .A1(n17005), .A2(n17661), .ZN(\DataMem/N2109 ) );
  AOI22_X1 U11623 ( .A1(n16823), .A2(\DataMem/Mem[7][7] ), .B1(n16824), .B2(
        \DataMem/Mem[6][7] ), .ZN(n16941) );
  AOI22_X1 U11622 ( .A1(n17531), .A2(\DataMem/Mem[5][7] ), .B1(n16822), .B2(
        \DataMem/Mem[4][7] ), .ZN(n16942) );
  AOI22_X1 U11621 ( .A1(n16819), .A2(\DataMem/Mem[3][7] ), .B1(n17653), .B2(
        \DataMem/Mem[2][7] ), .ZN(n16943) );
  AOI22_X1 U11620 ( .A1(n17124), .A2(\DataMem/Mem[1][7] ), .B1(n17125), .B2(
        \DataMem/Mem[0][7] ), .ZN(n16944) );
  NOR2_X1 U11618 ( .A1(n17155), .A2(n16940), .ZN(\DataMem/N2182 ) );
  NOR2_X1 U11957 ( .A1(n17004), .A2(n17650), .ZN(\DataMem/N1663 ) );
  NOR2_X1 U11692 ( .A1(n17006), .A2(n17661), .ZN(\DataMem/N2107 ) );
  NOR2_X1 U11898 ( .A1(n17004), .A2(n17651), .ZN(\DataMem/N1727 ) );
  NOR2_X1 U11726 ( .A1(n17006), .A2(n17658), .ZN(\DataMem/N2043 ) );
  NOR2_X1 U11761 ( .A1(n17006), .A2(n17657), .ZN(\DataMem/N1979 ) );
  NOR2_X1 U11863 ( .A1(n17004), .A2(n17654), .ZN(\DataMem/N1791 ) );
  NOR2_X1 U11796 ( .A1(n17006), .A2(n17656), .ZN(\DataMem/N1915 ) );
  NOR2_X1 U11830 ( .A1(n17006), .A2(n17655), .ZN(\DataMem/N1851 ) );
  NOR2_X1 U11828 ( .A1(n17004), .A2(n17655), .ZN(\DataMem/N1855 ) );
  NOR2_X1 U11865 ( .A1(n17006), .A2(n17654), .ZN(\DataMem/N1787 ) );
  NOR2_X1 U11900 ( .A1(n17006), .A2(n17651), .ZN(\DataMem/N1723 ) );
  NOR2_X1 U11794 ( .A1(n17004), .A2(n17656), .ZN(\DataMem/N1919 ) );
  NOR2_X1 U11961 ( .A1(n17006), .A2(n17650), .ZN(\DataMem/N1659 ) );
  AOI22_X1 U11635 ( .A1(n16823), .A2(\DataMem/Mem[7][5] ), .B1(n17530), .B2(
        \DataMem/Mem[6][5] ), .ZN(n16951) );
  AOI22_X1 U11634 ( .A1(n17531), .A2(\DataMem/Mem[5][5] ), .B1(n16822), .B2(
        \DataMem/Mem[4][5] ), .ZN(n16952) );
  AOI22_X1 U11633 ( .A1(n17122), .A2(\DataMem/Mem[3][5] ), .B1(n17652), .B2(
        \DataMem/Mem[2][5] ), .ZN(n16953) );
  AOI22_X1 U11632 ( .A1(n17124), .A2(\DataMem/Mem[1][5] ), .B1(n16818), .B2(
        \DataMem/Mem[0][5] ), .ZN(n16954) );
  NOR2_X1 U11630 ( .A1(n17155), .A2(n16950), .ZN(\DataMem/N2176 ) );
  NOR2_X1 U11824 ( .A1(n17000), .A2(n16594), .ZN(\DataMem/N1863 ) );
  NOR2_X1 U11790 ( .A1(n17000), .A2(n16593), .ZN(\DataMem/N1927 ) );
  NOR2_X1 U11755 ( .A1(n17000), .A2(n16592), .ZN(\DataMem/N1991 ) );
  NOR2_X1 U11720 ( .A1(n17000), .A2(n16591), .ZN(\DataMem/N2055 ) );
  NOR2_X1 U11686 ( .A1(n17000), .A2(n16590), .ZN(\DataMem/N2119 ) );
  AOI22_X1 U11611 ( .A1(n17660), .A2(\DataMem/Mem[7][9] ), .B1(n16824), .B2(
        \DataMem/Mem[6][9] ), .ZN(n16931) );
  AOI22_X1 U11610 ( .A1(n16821), .A2(\DataMem/Mem[5][9] ), .B1(n16822), .B2(
        \DataMem/Mem[4][9] ), .ZN(n16932) );
  AOI22_X1 U11609 ( .A1(n17122), .A2(\DataMem/Mem[3][9] ), .B1(n17653), .B2(
        \DataMem/Mem[2][9] ), .ZN(n16933) );
  AOI22_X1 U11608 ( .A1(n17124), .A2(\DataMem/Mem[1][9] ), .B1(n16818), .B2(
        \DataMem/Mem[0][9] ), .ZN(n16934) );
  NOR2_X1 U11606 ( .A1(n17155), .A2(n16930), .ZN(\DataMem/N2188 ) );
  NOR2_X1 U11953 ( .A1(n17002), .A2(n16597), .ZN(\DataMem/N1667 ) );
  NOR2_X1 U11896 ( .A1(n17002), .A2(n16596), .ZN(\DataMem/N1731 ) );
  NOR2_X1 U11861 ( .A1(n17002), .A2(n16595), .ZN(\DataMem/N1795 ) );
  NOR2_X1 U11826 ( .A1(n17002), .A2(n16594), .ZN(\DataMem/N1859 ) );
  NOR2_X1 U11792 ( .A1(n17002), .A2(n16593), .ZN(\DataMem/N1923 ) );
  NOR2_X1 U11757 ( .A1(n17002), .A2(n16592), .ZN(\DataMem/N1987 ) );
  NOR2_X1 U11722 ( .A1(n17002), .A2(n16591), .ZN(\DataMem/N2051 ) );
  NOR2_X1 U11688 ( .A1(n17002), .A2(n16590), .ZN(\DataMem/N2115 ) );
  NOR2_X1 U11969 ( .A1(n17010), .A2(n17650), .ZN(\DataMem/N1651 ) );
  AOI22_X1 U11659 ( .A1(n17659), .A2(\DataMem/Mem[7][1] ), .B1(n17530), .B2(
        \DataMem/Mem[6][1] ), .ZN(n16971) );
  AOI22_X1 U11658 ( .A1(n17531), .A2(\DataMem/Mem[5][1] ), .B1(n16822), .B2(
        \DataMem/Mem[4][1] ), .ZN(n16972) );
  AOI22_X1 U11657 ( .A1(n17122), .A2(\DataMem/Mem[3][1] ), .B1(n17653), .B2(
        \DataMem/Mem[2][1] ), .ZN(n16973) );
  AOI22_X1 U11656 ( .A1(n17124), .A2(\DataMem/Mem[1][1] ), .B1(n17125), .B2(
        \DataMem/Mem[0][1] ), .ZN(n16974) );
  NOR2_X1 U11654 ( .A1(n17155), .A2(n16970), .ZN(\DataMem/N2164 ) );
  NOR2_X1 U11959 ( .A1(n17005), .A2(n17650), .ZN(\DataMem/N1661 ) );
  AOI22_X1 U11629 ( .A1(n16823), .A2(\DataMem/Mem[7][6] ), .B1(n17530), .B2(
        \DataMem/Mem[6][6] ), .ZN(n16946) );
  AOI22_X1 U11628 ( .A1(n17531), .A2(\DataMem/Mem[5][6] ), .B1(n16822), .B2(
        \DataMem/Mem[4][6] ), .ZN(n16947) );
  AOI22_X1 U11627 ( .A1(n16819), .A2(\DataMem/Mem[3][6] ), .B1(n17652), .B2(
        \DataMem/Mem[2][6] ), .ZN(n16948) );
  AOI22_X1 U11626 ( .A1(n17124), .A2(\DataMem/Mem[1][6] ), .B1(n17125), .B2(
        \DataMem/Mem[0][6] ), .ZN(n16949) );
  NOR2_X1 U11624 ( .A1(n17155), .A2(n16945), .ZN(\DataMem/N2179 ) );
  NOR2_X1 U11690 ( .A1(n17004), .A2(n17661), .ZN(\DataMem/N2111 ) );
  NOR2_X1 U11771 ( .A1(n16981), .A2(n17656), .ZN(\DataMem/N1965 ) );
  NOR2_X1 U11897 ( .A1(n17003), .A2(n16596), .ZN(\DataMem/N1729 ) );
  NOR2_X1 U11736 ( .A1(n16981), .A2(n17657), .ZN(\DataMem/N2029 ) );
  NOR2_X1 U11701 ( .A1(n16981), .A2(n17658), .ZN(\DataMem/N2093 ) );
  NOR2_X1 U11667 ( .A1(n16981), .A2(n17661), .ZN(\DataMem/N2157 ) );
  NOR2_X1 U11955 ( .A1(n17003), .A2(n16597), .ZN(\DataMem/N1665 ) );
  AOI22_X1 U11491 ( .A1(n16823), .A2(\DataMem/Mem[7][29] ), .B1(n16824), .B2(
        \DataMem/Mem[6][29] ), .ZN(n16831) );
  AOI22_X1 U11490 ( .A1(n17531), .A2(\DataMem/Mem[5][29] ), .B1(n16822), .B2(
        \DataMem/Mem[4][29] ), .ZN(n16832) );
  AOI22_X1 U11489 ( .A1(n17122), .A2(\DataMem/Mem[3][29] ), .B1(n17653), .B2(
        \DataMem/Mem[2][29] ), .ZN(n16833) );
  AOI22_X1 U11488 ( .A1(n16817), .A2(\DataMem/Mem[1][29] ), .B1(n17125), .B2(
        \DataMem/Mem[0][29] ), .ZN(n16834) );
  NOR2_X1 U11486 ( .A1(n17155), .A2(n16830), .ZN(\DataMem/N2248 ) );
  NOR2_X1 U11913 ( .A1(n16982), .A2(n17650), .ZN(\DataMem/N1707 ) );
  AOI22_X1 U11617 ( .A1(n17659), .A2(\DataMem/Mem[7][8] ), .B1(n16824), .B2(
        \DataMem/Mem[6][8] ), .ZN(n16936) );
  AOI22_X1 U11616 ( .A1(n17531), .A2(\DataMem/Mem[5][8] ), .B1(n16822), .B2(
        \DataMem/Mem[4][8] ), .ZN(n16937) );
  AOI22_X1 U11615 ( .A1(n17122), .A2(\DataMem/Mem[3][8] ), .B1(n17653), .B2(
        \DataMem/Mem[2][8] ), .ZN(n16938) );
  AOI22_X1 U11614 ( .A1(n16817), .A2(\DataMem/Mem[1][8] ), .B1(n16818), .B2(
        \DataMem/Mem[0][8] ), .ZN(n16939) );
  NOR2_X1 U11612 ( .A1(n17155), .A2(n16935), .ZN(\DataMem/N2185 ) );
  NOR2_X1 U11876 ( .A1(n16982), .A2(n17651), .ZN(\DataMem/N1771 ) );
  NOR2_X1 U11841 ( .A1(n16982), .A2(n17654), .ZN(\DataMem/N1835 ) );
  NOR2_X1 U11806 ( .A1(n16982), .A2(n17655), .ZN(\DataMem/N1899 ) );
  NOR2_X1 U11772 ( .A1(n16982), .A2(n17656), .ZN(\DataMem/N1963 ) );
  NOR2_X1 U11697 ( .A1(n17011), .A2(n17661), .ZN(\DataMem/N2097 ) );
  NOR2_X1 U11737 ( .A1(n16982), .A2(n17657), .ZN(\DataMem/N2027 ) );
  NOR2_X1 U11702 ( .A1(n16982), .A2(n17658), .ZN(\DataMem/N2091 ) );
  NOR2_X1 U11668 ( .A1(n16982), .A2(n17661), .ZN(\DataMem/N2155 ) );
  NOR2_X1 U11731 ( .A1(n17011), .A2(n17658), .ZN(\DataMem/N2033 ) );
  AOI22_X1 U11503 ( .A1(n16823), .A2(\DataMem/Mem[7][27] ), .B1(n17530), .B2(
        \DataMem/Mem[6][27] ), .ZN(n16841) );
  AOI22_X1 U11502 ( .A1(n17531), .A2(\DataMem/Mem[5][27] ), .B1(n16822), .B2(
        \DataMem/Mem[4][27] ), .ZN(n16842) );
  AOI22_X1 U11501 ( .A1(n17122), .A2(\DataMem/Mem[3][27] ), .B1(n17653), .B2(
        \DataMem/Mem[2][27] ), .ZN(n16843) );
  AOI22_X1 U11500 ( .A1(n17124), .A2(\DataMem/Mem[1][27] ), .B1(n17125), .B2(
        \DataMem/Mem[0][27] ), .ZN(n16844) );
  NOR2_X1 U11498 ( .A1(n17155), .A2(n16840), .ZN(\DataMem/N2242 ) );
  AOI22_X1 U11918 ( .A1(\pipeline/Forward_sw1_mux ), .A2(
        \pipeline/data_to_RF_from_WB[27] ), .B1(n13793), .B2(n17743), .ZN(
        n16984) );
  NOR2_X1 U11917 ( .A1(n16984), .A2(n17650), .ZN(\DataMem/N1703 ) );
  NOR2_X1 U11878 ( .A1(n16984), .A2(n17651), .ZN(\DataMem/N1767 ) );
  NOR2_X1 U11766 ( .A1(n17011), .A2(n17657), .ZN(\DataMem/N1969 ) );
  NOR2_X1 U11843 ( .A1(n16984), .A2(n17654), .ZN(\DataMem/N1831 ) );
  NOR2_X1 U11808 ( .A1(n16984), .A2(n17655), .ZN(\DataMem/N1895 ) );
  NOR2_X1 U11774 ( .A1(n16984), .A2(n17656), .ZN(\DataMem/N1959 ) );
  NOR2_X1 U11801 ( .A1(n17011), .A2(n17656), .ZN(\DataMem/N1905 ) );
  NOR2_X1 U11739 ( .A1(n16984), .A2(n17657), .ZN(\DataMem/N2023 ) );
  NOR2_X1 U11672 ( .A1(n16986), .A2(n16590), .ZN(\DataMem/N2147 ) );
  NOR2_X1 U11704 ( .A1(n16984), .A2(n17658), .ZN(\DataMem/N2087 ) );
  NOR2_X1 U11670 ( .A1(n16984), .A2(n17661), .ZN(\DataMem/N2151 ) );
  NOR2_X1 U11835 ( .A1(n17011), .A2(n17655), .ZN(\DataMem/N1841 ) );
  AOI22_X1 U11509 ( .A1(n17660), .A2(\DataMem/Mem[7][26] ), .B1(n17530), .B2(
        \DataMem/Mem[6][26] ), .ZN(n16846) );
  AOI22_X1 U11508 ( .A1(n17531), .A2(\DataMem/Mem[5][26] ), .B1(n16822), .B2(
        \DataMem/Mem[4][26] ), .ZN(n16847) );
  AOI22_X1 U11507 ( .A1(n17122), .A2(\DataMem/Mem[3][26] ), .B1(n17652), .B2(
        \DataMem/Mem[2][26] ), .ZN(n16848) );
  AOI22_X1 U11506 ( .A1(n17124), .A2(\DataMem/Mem[1][26] ), .B1(n17125), .B2(
        \DataMem/Mem[0][26] ), .ZN(n16849) );
  NOR2_X1 U11504 ( .A1(n17155), .A2(n16845), .ZN(\DataMem/N2239 ) );
  AOI22_X1 U11920 ( .A1(\pipeline/Forward_sw1_mux ), .A2(
        \pipeline/data_to_RF_from_WB[26] ), .B1(n13794), .B2(n17380), .ZN(
        n16985) );
  NOR2_X1 U11919 ( .A1(n16985), .A2(n17650), .ZN(\DataMem/N1701 ) );
  NOR2_X1 U11870 ( .A1(n17011), .A2(n17654), .ZN(\DataMem/N1777 ) );
  NOR2_X1 U11879 ( .A1(n16985), .A2(n17651), .ZN(\DataMem/N1765 ) );
  NOR2_X1 U11844 ( .A1(n16985), .A2(n17654), .ZN(\DataMem/N1829 ) );
  NOR2_X1 U11809 ( .A1(n16985), .A2(n17655), .ZN(\DataMem/N1893 ) );
  NOR2_X1 U11905 ( .A1(n17011), .A2(n17651), .ZN(\DataMem/N1713 ) );
  NOR2_X1 U11775 ( .A1(n16985), .A2(n17656), .ZN(\DataMem/N1957 ) );
  NOR2_X1 U11740 ( .A1(n16985), .A2(n17657), .ZN(\DataMem/N2021 ) );
  NOR2_X1 U11705 ( .A1(n16985), .A2(n17658), .ZN(\DataMem/N2085 ) );
  NOR2_X1 U11971 ( .A1(n17011), .A2(n17650), .ZN(\DataMem/N1649 ) );
  NOR2_X1 U11671 ( .A1(n16985), .A2(n17661), .ZN(\DataMem/N2149 ) );
  AOI22_X1 U11665 ( .A1(n17659), .A2(\DataMem/Mem[7][0] ), .B1(n17530), .B2(
        \DataMem/Mem[6][0] ), .ZN(n16976) );
  AOI22_X1 U11664 ( .A1(n17531), .A2(\DataMem/Mem[5][0] ), .B1(n16822), .B2(
        \DataMem/Mem[4][0] ), .ZN(n16977) );
  AOI22_X1 U11663 ( .A1(n17122), .A2(\DataMem/Mem[3][0] ), .B1(n17652), .B2(
        \DataMem/Mem[2][0] ), .ZN(n16978) );
  AOI22_X1 U11662 ( .A1(n17124), .A2(\DataMem/Mem[1][0] ), .B1(n17125), .B2(
        \DataMem/Mem[0][0] ), .ZN(n16979) );
  NOR2_X1 U11660 ( .A1(n17155), .A2(n16975), .ZN(\DataMem/N2161 ) );
  AOI22_X1 U11515 ( .A1(n17660), .A2(\DataMem/Mem[7][25] ), .B1(n17530), .B2(
        \DataMem/Mem[6][25] ), .ZN(n16851) );
  AOI22_X1 U11514 ( .A1(n17531), .A2(\DataMem/Mem[5][25] ), .B1(n16822), .B2(
        \DataMem/Mem[4][25] ), .ZN(n16852) );
  AOI22_X1 U11513 ( .A1(n17122), .A2(\DataMem/Mem[3][25] ), .B1(n16820), .B2(
        \DataMem/Mem[2][25] ), .ZN(n16853) );
  AOI22_X1 U11512 ( .A1(n17124), .A2(\DataMem/Mem[1][25] ), .B1(n16818), .B2(
        \DataMem/Mem[0][25] ), .ZN(n16854) );
  NOR2_X1 U11510 ( .A1(n17155), .A2(n16850), .ZN(\DataMem/N2236 ) );
  NOR2_X1 U11921 ( .A1(n16986), .A2(n16597), .ZN(\DataMem/N1699 ) );
  NOR2_X1 U11880 ( .A1(n16986), .A2(n16596), .ZN(\DataMem/N1763 ) );
  AOI22_X1 U11910 ( .A1(\pipeline/Forward_sw1_mux ), .A2(
        \pipeline/data_to_RF_from_WB[31] ), .B1(n13783), .B2(n17380), .ZN(
        n16980) );
  NOR2_X1 U11700 ( .A1(n16980), .A2(n17658), .ZN(\DataMem/N2095 ) );
  NOR2_X1 U11845 ( .A1(n16986), .A2(n16595), .ZN(\DataMem/N1827 ) );
  NOR2_X1 U11810 ( .A1(n16986), .A2(n16594), .ZN(\DataMem/N1891 ) );
  NOR2_X1 U11735 ( .A1(n16980), .A2(n17657), .ZN(\DataMem/N2031 ) );
  NOR2_X1 U11776 ( .A1(n16986), .A2(n16593), .ZN(\DataMem/N1955 ) );
  NOR2_X1 U11741 ( .A1(n16986), .A2(n16592), .ZN(\DataMem/N2019 ) );
  NOR2_X1 U11706 ( .A1(n16986), .A2(n16591), .ZN(\DataMem/N2083 ) );
  NOR2_X1 U11770 ( .A1(n16980), .A2(n17656), .ZN(\DataMem/N1967 ) );
  NOR2_X1 U11915 ( .A1(n16983), .A2(n17650), .ZN(\DataMem/N1705 ) );
  NOR2_X1 U11877 ( .A1(n16983), .A2(n17651), .ZN(\DataMem/N1769 ) );
  NOR2_X1 U11673 ( .A1(n16987), .A2(n16590), .ZN(\DataMem/N2145 ) );
  NOR2_X1 U11842 ( .A1(n16983), .A2(n17654), .ZN(\DataMem/N1833 ) );
  NOR2_X1 U11807 ( .A1(n16983), .A2(n17655), .ZN(\DataMem/N1897 ) );
  NOR2_X1 U11773 ( .A1(n16983), .A2(n17656), .ZN(\DataMem/N1961 ) );
  NOR2_X1 U11707 ( .A1(n16987), .A2(n16591), .ZN(\DataMem/N2081 ) );
  NOR2_X1 U11738 ( .A1(n16983), .A2(n17657), .ZN(\DataMem/N2025 ) );
  NOR2_X1 U11703 ( .A1(n16983), .A2(n17658), .ZN(\DataMem/N2089 ) );
  NOR2_X1 U11742 ( .A1(n16987), .A2(n16592), .ZN(\DataMem/N2017 ) );
  NOR2_X1 U11669 ( .A1(n16983), .A2(n17661), .ZN(\DataMem/N2153 ) );
  AOI22_X1 U11581 ( .A1(n17659), .A2(\DataMem/Mem[7][14] ), .B1(n17530), .B2(
        \DataMem/Mem[6][14] ), .ZN(n16906) );
  AOI22_X1 U11580 ( .A1(n16821), .A2(\DataMem/Mem[5][14] ), .B1(n16822), .B2(
        \DataMem/Mem[4][14] ), .ZN(n16907) );
  AOI22_X1 U11579 ( .A1(n17122), .A2(\DataMem/Mem[3][14] ), .B1(n17653), .B2(
        \DataMem/Mem[2][14] ), .ZN(n16908) );
  AOI22_X1 U11578 ( .A1(n17124), .A2(\DataMem/Mem[1][14] ), .B1(n16818), .B2(
        \DataMem/Mem[0][14] ), .ZN(n16909) );
  NOR2_X1 U11576 ( .A1(n17155), .A2(n16905), .ZN(\DataMem/N2203 ) );
  NOR2_X1 U11943 ( .A1(n16997), .A2(n17650), .ZN(\DataMem/N1677 ) );
  NOR2_X1 U11891 ( .A1(n16997), .A2(n17651), .ZN(\DataMem/N1741 ) );
  NOR2_X1 U11777 ( .A1(n16987), .A2(n16593), .ZN(\DataMem/N1953 ) );
  NOR2_X1 U11856 ( .A1(n16997), .A2(n17654), .ZN(\DataMem/N1805 ) );
  NOR2_X1 U11821 ( .A1(n16997), .A2(n17655), .ZN(\DataMem/N1869 ) );
  NOR2_X1 U11787 ( .A1(n16997), .A2(n17656), .ZN(\DataMem/N1933 ) );
  NOR2_X1 U11811 ( .A1(n16987), .A2(n16594), .ZN(\DataMem/N1889 ) );
  NOR2_X1 U11752 ( .A1(n16997), .A2(n17657), .ZN(\DataMem/N1997 ) );
  NOR2_X1 U11717 ( .A1(n16997), .A2(n17658), .ZN(\DataMem/N2061 ) );
  NOR2_X1 U11846 ( .A1(n16987), .A2(n16595), .ZN(\DataMem/N1825 ) );
  NOR2_X1 U11683 ( .A1(n16997), .A2(n17661), .ZN(\DataMem/N2125 ) );
  AOI22_X1 U11575 ( .A1(n17659), .A2(\DataMem/Mem[7][15] ), .B1(n16824), .B2(
        \DataMem/Mem[6][15] ), .ZN(n16901) );
  AOI22_X1 U11574 ( .A1(n16821), .A2(\DataMem/Mem[5][15] ), .B1(n16822), .B2(
        \DataMem/Mem[4][15] ), .ZN(n16902) );
  AOI22_X1 U11573 ( .A1(n17122), .A2(\DataMem/Mem[3][15] ), .B1(n17653), .B2(
        \DataMem/Mem[2][15] ), .ZN(n16903) );
  AOI22_X1 U11572 ( .A1(n16817), .A2(\DataMem/Mem[1][15] ), .B1(n17125), .B2(
        \DataMem/Mem[0][15] ), .ZN(n16904) );
  NOR2_X1 U11570 ( .A1(n12766), .A2(n16900), .ZN(\DataMem/N2206 ) );
  NOR2_X1 U11881 ( .A1(n16987), .A2(n16596), .ZN(\DataMem/N1761 ) );
  NOR2_X1 U11941 ( .A1(n16996), .A2(n17650), .ZN(\DataMem/N1679 ) );
  NOR2_X1 U11890 ( .A1(n16996), .A2(n17651), .ZN(\DataMem/N1743 ) );
  NOR2_X1 U11855 ( .A1(n16996), .A2(n17654), .ZN(\DataMem/N1807 ) );
  NOR2_X1 U11923 ( .A1(n16987), .A2(n16597), .ZN(\DataMem/N1697 ) );
  NOR2_X1 U11820 ( .A1(n16996), .A2(n17655), .ZN(\DataMem/N1871 ) );
  AOI22_X1 U11521 ( .A1(n17660), .A2(\DataMem/Mem[7][24] ), .B1(n17530), .B2(
        \DataMem/Mem[6][24] ), .ZN(n16856) );
  AOI22_X1 U11520 ( .A1(n17531), .A2(\DataMem/Mem[5][24] ), .B1(n16822), .B2(
        \DataMem/Mem[4][24] ), .ZN(n16857) );
  AOI22_X1 U11519 ( .A1(n16819), .A2(\DataMem/Mem[3][24] ), .B1(n16820), .B2(
        \DataMem/Mem[2][24] ), .ZN(n16858) );
  AOI22_X1 U11518 ( .A1(n16817), .A2(\DataMem/Mem[1][24] ), .B1(n16818), .B2(
        \DataMem/Mem[0][24] ), .ZN(n16859) );
  NOR2_X1 U11516 ( .A1(n17155), .A2(n16855), .ZN(\DataMem/N2233 ) );
  NOR2_X1 U11786 ( .A1(n16996), .A2(n17656), .ZN(\DataMem/N1935 ) );
  NOR2_X1 U11751 ( .A1(n16996), .A2(n17657), .ZN(\DataMem/N1999 ) );
  NOR2_X1 U11716 ( .A1(n16996), .A2(n17658), .ZN(\DataMem/N2063 ) );
  NOR2_X1 U11689 ( .A1(n17003), .A2(n16590), .ZN(\DataMem/N2113 ) );
  NOR2_X1 U11682 ( .A1(n16996), .A2(n17661), .ZN(\DataMem/N2127 ) );
  AOI22_X1 U11587 ( .A1(n17659), .A2(\DataMem/Mem[7][13] ), .B1(n16824), .B2(
        \DataMem/Mem[6][13] ), .ZN(n16911) );
  AOI22_X1 U11586 ( .A1(n16821), .A2(\DataMem/Mem[5][13] ), .B1(n16822), .B2(
        \DataMem/Mem[4][13] ), .ZN(n16912) );
  AOI22_X1 U11585 ( .A1(n17122), .A2(\DataMem/Mem[3][13] ), .B1(n17653), .B2(
        \DataMem/Mem[2][13] ), .ZN(n16913) );
  AOI22_X1 U11584 ( .A1(n16817), .A2(\DataMem/Mem[1][13] ), .B1(n17125), .B2(
        \DataMem/Mem[0][13] ), .ZN(n16914) );
  NOR2_X1 U11582 ( .A1(n12766), .A2(n16910), .ZN(\DataMem/N2200 ) );
  AOI22_X1 U11946 ( .A1(\pipeline/Forward_sw1_mux ), .A2(
        \pipeline/data_to_RF_from_WB[13] ), .B1(n13790), .B2(n17380), .ZN(
        n16998) );
  NOR2_X1 U11945 ( .A1(n16998), .A2(n17650), .ZN(\DataMem/N1675 ) );
  NOR2_X1 U11723 ( .A1(n17003), .A2(n16591), .ZN(\DataMem/N2049 ) );
  NOR2_X1 U11892 ( .A1(n16998), .A2(n17651), .ZN(\DataMem/N1739 ) );
  NOR2_X1 U11857 ( .A1(n16998), .A2(n17654), .ZN(\DataMem/N1803 ) );
  NOR2_X1 U11758 ( .A1(n17003), .A2(n16592), .ZN(\DataMem/N1985 ) );
  NOR2_X1 U11822 ( .A1(n16998), .A2(n17655), .ZN(\DataMem/N1867 ) );
  NOR2_X1 U11788 ( .A1(n16998), .A2(n17656), .ZN(\DataMem/N1931 ) );
  NOR2_X1 U11753 ( .A1(n16998), .A2(n17657), .ZN(\DataMem/N1995 ) );
  NOR2_X1 U11793 ( .A1(n17003), .A2(n16593), .ZN(\DataMem/N1921 ) );
  NOR2_X1 U11718 ( .A1(n16998), .A2(n17658), .ZN(\DataMem/N2059 ) );
  NOR2_X1 U11684 ( .A1(n16998), .A2(n17661), .ZN(\DataMem/N2123 ) );
  NOR2_X1 U11827 ( .A1(n17003), .A2(n16594), .ZN(\DataMem/N1857 ) );
  AOI22_X1 U11485 ( .A1(n17659), .A2(\DataMem/Mem[7][30] ), .B1(n16824), .B2(
        \DataMem/Mem[6][30] ), .ZN(n16826) );
  AOI22_X1 U11484 ( .A1(n17531), .A2(\DataMem/Mem[5][30] ), .B1(n16822), .B2(
        \DataMem/Mem[4][30] ), .ZN(n16827) );
  AOI22_X1 U11483 ( .A1(n17122), .A2(\DataMem/Mem[3][30] ), .B1(n17653), .B2(
        \DataMem/Mem[2][30] ), .ZN(n16828) );
  AOI22_X1 U11482 ( .A1(n17124), .A2(\DataMem/Mem[1][30] ), .B1(n16818), .B2(
        \DataMem/Mem[0][30] ), .ZN(n16829) );
  NOR2_X1 U11480 ( .A1(n17155), .A2(n16825), .ZN(\DataMem/N2251 ) );
  NOR2_X1 U11911 ( .A1(n16981), .A2(n17650), .ZN(\DataMem/N1709 ) );
  NOR2_X1 U11875 ( .A1(n16981), .A2(n17651), .ZN(\DataMem/N1773 ) );
  NOR2_X1 U11840 ( .A1(n16981), .A2(n17654), .ZN(\DataMem/N1837 ) );
  NOR2_X1 U11862 ( .A1(n17003), .A2(n16595), .ZN(\DataMem/N1793 ) );
  NOR2_X1 U11805 ( .A1(n16981), .A2(n17655), .ZN(\DataMem/N1901 ) );
  NOR2_X1 U11724 ( .A1(n17004), .A2(n17658), .ZN(\DataMem/N2047 ) );
  AOI22_X1 U11497 ( .A1(n16823), .A2(\DataMem/Mem[7][28] ), .B1(n17530), .B2(
        \DataMem/Mem[6][28] ), .ZN(n16836) );
  AOI22_X1 U11496 ( .A1(n17531), .A2(\DataMem/Mem[5][28] ), .B1(n16822), .B2(
        \DataMem/Mem[4][28] ), .ZN(n16837) );
  AOI22_X1 U11495 ( .A1(n17122), .A2(\DataMem/Mem[3][28] ), .B1(n17653), .B2(
        \DataMem/Mem[2][28] ), .ZN(n16838) );
  AOI22_X1 U11494 ( .A1(n17124), .A2(\DataMem/Mem[1][28] ), .B1(n17125), .B2(
        \DataMem/Mem[0][28] ), .ZN(n16839) );
  NOR2_X1 U11492 ( .A1(n12766), .A2(n16835), .ZN(\DataMem/N2245 ) );
  NOR2_X1 U11710 ( .A1(n16990), .A2(n16591), .ZN(\DataMem/N2075 ) );
  NOR2_X1 U11818 ( .A1(n16994), .A2(n16594), .ZN(\DataMem/N1875 ) );
  NOR2_X1 U11676 ( .A1(n16990), .A2(n16590), .ZN(\DataMem/N2139 ) );
  AOI22_X1 U11545 ( .A1(n17660), .A2(\DataMem/Mem[7][20] ), .B1(n17530), .B2(
        \DataMem/Mem[6][20] ), .ZN(n16876) );
  AOI22_X1 U11544 ( .A1(n16821), .A2(\DataMem/Mem[5][20] ), .B1(n16822), .B2(
        \DataMem/Mem[4][20] ), .ZN(n16877) );
  AOI22_X1 U11543 ( .A1(n16819), .A2(\DataMem/Mem[3][20] ), .B1(n17653), .B2(
        \DataMem/Mem[2][20] ), .ZN(n16878) );
  AOI22_X1 U11542 ( .A1(n17124), .A2(\DataMem/Mem[1][20] ), .B1(n17125), .B2(
        \DataMem/Mem[0][20] ), .ZN(n16879) );
  NOR2_X1 U11540 ( .A1(n17155), .A2(n16875), .ZN(\DataMem/N2221 ) );
  NOR2_X1 U11931 ( .A1(n16991), .A2(n16597), .ZN(\DataMem/N1689 ) );
  NOR2_X1 U11885 ( .A1(n16991), .A2(n16596), .ZN(\DataMem/N1753 ) );
  NOR2_X1 U11850 ( .A1(n16991), .A2(n16595), .ZN(\DataMem/N1817 ) );
  NOR2_X1 U11815 ( .A1(n16991), .A2(n16594), .ZN(\DataMem/N1881 ) );
  NOR2_X1 U11781 ( .A1(n16991), .A2(n16593), .ZN(\DataMem/N1945 ) );
  NOR2_X1 U11853 ( .A1(n16994), .A2(n16595), .ZN(\DataMem/N1811 ) );
  NOR2_X1 U11746 ( .A1(n16991), .A2(n16592), .ZN(\DataMem/N2009 ) );
  NOR2_X1 U11711 ( .A1(n16991), .A2(n16591), .ZN(\DataMem/N2073 ) );
  NOR2_X1 U11677 ( .A1(n16991), .A2(n16590), .ZN(\DataMem/N2137 ) );
  AOI22_X1 U11551 ( .A1(n17659), .A2(\DataMem/Mem[7][19] ), .B1(n16824), .B2(
        \DataMem/Mem[6][19] ), .ZN(n16881) );
  AOI22_X1 U11550 ( .A1(n16821), .A2(\DataMem/Mem[5][19] ), .B1(n16822), .B2(
        \DataMem/Mem[4][19] ), .ZN(n16882) );
  AOI22_X1 U11549 ( .A1(n17122), .A2(\DataMem/Mem[3][19] ), .B1(n16820), .B2(
        \DataMem/Mem[2][19] ), .ZN(n16883) );
  AOI22_X1 U11548 ( .A1(n17124), .A2(\DataMem/Mem[1][19] ), .B1(n16818), .B2(
        \DataMem/Mem[0][19] ), .ZN(n16884) );
  NOR2_X1 U11546 ( .A1(n17155), .A2(n16880), .ZN(\DataMem/N2218 ) );
  NOR2_X1 U11888 ( .A1(n16994), .A2(n16596), .ZN(\DataMem/N1747 ) );
  AOI22_X1 U11934 ( .A1(\pipeline/Forward_sw1_mux ), .A2(
        \pipeline/data_to_RF_from_WB[19] ), .B1(n13800), .B2(n17380), .ZN(
        n16992) );
  NOR2_X1 U11933 ( .A1(n16992), .A2(n16597), .ZN(\DataMem/N1687 ) );
  NOR2_X1 U11886 ( .A1(n16992), .A2(n16596), .ZN(\DataMem/N1751 ) );
  AOI22_X1 U11936 ( .A1(\pipeline/Forward_sw1_mux ), .A2(
        \pipeline/data_to_RF_from_WB[18] ), .B1(n13801), .B2(n17380), .ZN(
        n16993) );
  NOR2_X1 U11713 ( .A1(n16993), .A2(n16591), .ZN(\DataMem/N2069 ) );
  NOR2_X1 U11851 ( .A1(n16992), .A2(n16595), .ZN(\DataMem/N1815 ) );
  NOR2_X1 U11816 ( .A1(n16992), .A2(n16594), .ZN(\DataMem/N1879 ) );
  NOR2_X1 U11937 ( .A1(n16994), .A2(n16597), .ZN(\DataMem/N1683 ) );
  NOR2_X1 U11782 ( .A1(n16992), .A2(n16593), .ZN(\DataMem/N1943 ) );
  AOI22_X1 U11563 ( .A1(n17660), .A2(\DataMem/Mem[7][17] ), .B1(n16824), .B2(
        \DataMem/Mem[6][17] ), .ZN(n16891) );
  AOI22_X1 U11562 ( .A1(n16821), .A2(\DataMem/Mem[5][17] ), .B1(n16822), .B2(
        \DataMem/Mem[4][17] ), .ZN(n16892) );
  AOI22_X1 U11561 ( .A1(n17122), .A2(\DataMem/Mem[3][17] ), .B1(n16820), .B2(
        \DataMem/Mem[2][17] ), .ZN(n16893) );
  AOI22_X1 U11560 ( .A1(n17124), .A2(\DataMem/Mem[1][17] ), .B1(n17125), .B2(
        \DataMem/Mem[0][17] ), .ZN(n16894) );
  NOR2_X1 U11558 ( .A1(n17155), .A2(n16890), .ZN(\DataMem/N2212 ) );
  NOR2_X1 U11747 ( .A1(n16992), .A2(n16592), .ZN(\DataMem/N2007 ) );
  NAND4_X1 U8521 ( .A1(n14116), .A2(n14117), .A3(n14113), .A4(n14100), .ZN(
        n14121) );
  NOR2_X1 U8520 ( .A1(n14120), .A2(n14121), .ZN(n14096) );
  NOR4_X1 U8508 ( .A1(n14096), .A2(n14097), .A3(n14098), .A4(n14099), .ZN(
        n14095) );
  AOI22_X1 U8519 ( .A1(\pipeline/stageD/offset_jump_sign_ext [21]), .A2(n14116), .B1(\pipeline/stageD/offset_jump_sign_ext [22]), .B2(n14117), .ZN(n14119) );
  OAI221_X1 U8518 ( .B1(\pipeline/stageD/offset_jump_sign_ext [21]), .B2(
        n14116), .C1(\pipeline/stageD/offset_jump_sign_ext [22]), .C2(n14117), 
        .A(n14119), .ZN(n14087) );
  NAND2_X1 U8526 ( .A1(n14123), .A2(n17704), .ZN(n13983) );
  NOR2_X1 U8527 ( .A1(n17449), .A2(n14122), .ZN(n14093) );
  AOI22_X1 U8507 ( .A1(n14091), .A2(n14092), .B1(n14093), .B2(n14094), .ZN(
        n14088) );
  NOR2_X1 U8524 ( .A1(n14091), .A2(n14122), .ZN(n14090) );
  OAI211_X1 U8506 ( .C1(n14086), .C2(n14087), .A(n14088), .B(n14089), .ZN(
        \pipeline/cu_hazard/N40 ) );
  NOR2_X1 U11712 ( .A1(n16992), .A2(n16591), .ZN(\DataMem/N2071 ) );
  OAI21_X1 U8467 ( .B1(n14031), .B2(n14032), .A(n14033), .ZN(n14013) );
  NAND2_X1 U8491 ( .A1(n14005), .A2(n13990), .ZN(n14030) );
  NOR3_X1 U8465 ( .A1(n14027), .A2(n14015), .A3(n14007), .ZN(n14026) );
  NAND4_X1 U8464 ( .A1(n14025), .A2(n14013), .A3(n14002), .A4(n14026), .ZN(
        \pipeline/cu_pipeline/N105 ) );
  NOR2_X1 U11678 ( .A1(n16992), .A2(n16590), .ZN(\DataMem/N2135 ) );
  NOR2_X1 U8488 ( .A1(n17313), .A2(n14047), .ZN(n14000) );
  OAI221_X1 U8452 ( .B1(n13999), .B2(n14000), .C1(n13999), .C2(n14001), .A(
        n17704), .ZN(n13985) );
  NOR2_X1 U8451 ( .A1(n13281), .A2(n13998), .ZN(n13994) );
  NOR3_X1 U8469 ( .A1(n17347), .A2(n17409), .A3(n17313), .ZN(n13995) );
  OAI21_X1 U8450 ( .B1(n13281), .B2(n13997), .A(n13983), .ZN(n13996) );
  AOI221_X1 U8449 ( .B1(n13993), .B2(n13994), .C1(n13995), .C2(n13994), .A(
        n13996), .ZN(n13986) );
  NOR2_X1 U8448 ( .A1(n13281), .A2(n13984), .ZN(n13992) );
  OAI221_X1 U8447 ( .B1(n13989), .B2(n13990), .C1(n13989), .C2(n17076), .A(
        n13992), .ZN(n13987) );
  NAND4_X1 U8446 ( .A1(n13985), .A2(n13986), .A3(n13987), .A4(n13988), .ZN(
        \pipeline/cu_pipeline/N110 ) );
  AOI22_X1 U11557 ( .A1(n17659), .A2(\DataMem/Mem[7][18] ), .B1(n16824), .B2(
        \DataMem/Mem[6][18] ), .ZN(n16886) );
  AOI22_X1 U11556 ( .A1(n16821), .A2(\DataMem/Mem[5][18] ), .B1(n16822), .B2(
        \DataMem/Mem[4][18] ), .ZN(n16887) );
  AOI22_X1 U11555 ( .A1(n16819), .A2(\DataMem/Mem[3][18] ), .B1(n17653), .B2(
        \DataMem/Mem[2][18] ), .ZN(n16888) );
  AOI22_X1 U11554 ( .A1(n16817), .A2(\DataMem/Mem[1][18] ), .B1(n17125), .B2(
        \DataMem/Mem[0][18] ), .ZN(n16889) );
  NOR2_X1 U11552 ( .A1(n12766), .A2(n16885), .ZN(\DataMem/N2215 ) );
  NAND2_X1 U8442 ( .A1(n13980), .A2(n13981), .ZN(\pipeline/cu_pipeline/N88 )
         );
  NOR2_X1 U11935 ( .A1(n16993), .A2(n16597), .ZN(\DataMem/N1685 ) );
  NOR2_X1 U8490 ( .A1(n14047), .A2(n14058), .ZN(n14068) );
  OAI211_X1 U8487 ( .C1(n14012), .C2(n14024), .A(n14029), .B(n14070), .ZN(
        n14069) );
  NOR2_X1 U8486 ( .A1(n14068), .A2(n14069), .ZN(n14053) );
  OAI211_X1 U8475 ( .C1(n17406), .C2(n14030), .A(n14053), .B(n14041), .ZN(
        \pipeline/cu_pipeline/N102 ) );
  NOR2_X1 U11887 ( .A1(n16993), .A2(n16596), .ZN(\DataMem/N1749 ) );
  NOR2_X1 U11679 ( .A1(n16993), .A2(n16590), .ZN(\DataMem/N2133 ) );
  OAI22_X1 U8501 ( .A1(n13993), .A2(n17348), .B1(n14084), .B2(n17532), .ZN(
        n14083) );
  AOI211_X1 U8500 ( .C1(\pipeline/stageD/offset_to_jump_temp [10]), .C2(
        \pipeline/cu_pipeline/N89 ), .A(n14009), .B(n14083), .ZN(n14073) );
  AOI221_X1 U8499 ( .B1(\pipeline/inst_IFID_DEC[27] ), .B2(
        \pipeline/inst_IFID_DEC[26] ), .C1(n17313), .C2(n13993), .A(
        \pipeline/inst_IFID_DEC[29] ), .ZN(n14075) );
  OAI21_X1 U8498 ( .B1(\pipeline/stageD/offset_to_jump_temp [9]), .B2(
        \pipeline/stageD/offset_to_jump_temp [8]), .A(
        \pipeline/cu_pipeline/N89 ), .ZN(n14082) );
  OAI211_X1 U8497 ( .C1(\pipeline/inst_IFID_DEC[29] ), .C2(n17348), .A(n14082), 
        .B(n14058), .ZN(n14076) );
  AOI21_X1 U8495 ( .B1(n17361), .B2(n17412), .A(n13984), .ZN(n14077) );
  AOI21_X1 U8494 ( .B1(\pipeline/stageD/offset_to_jump_temp [5]), .B2(n17410), 
        .A(n13984), .ZN(n14078) );
  NOR4_X1 U8493 ( .A1(n14075), .A2(n14076), .A3(n14077), .A4(n14078), .ZN(
        n14074) );
  NAND4_X1 U8492 ( .A1(n14071), .A2(n14072), .A3(n14073), .A4(n14074), .ZN(
        \pipeline/cu_pipeline/N101 ) );
  NOR2_X1 U11852 ( .A1(n16993), .A2(n16595), .ZN(\DataMem/N1813 ) );
  AOI21_X1 U8463 ( .B1(n14023), .B2(n14024), .A(n14012), .ZN(n14010) );
  NAND4_X1 U8461 ( .A1(n14018), .A2(n14019), .A3(n14020), .A4(n14021), .ZN(
        n14017) );
  NOR4_X1 U8460 ( .A1(n14015), .A2(n14016), .A3(n14010), .A4(n14017), .ZN(
        n14014) );
  OAI211_X1 U8459 ( .C1(n14006), .C2(n14012), .A(n14013), .B(n14014), .ZN(
        \pipeline/cu_pipeline/N106 ) );
  OAI211_X1 U8468 ( .C1(n14023), .C2(n14012), .A(n14034), .B(n14035), .ZN(
        \pipeline/cu_pipeline/N104 ) );
  NOR2_X1 U11817 ( .A1(n16993), .A2(n16594), .ZN(\DataMem/N1877 ) );
  OAI21_X1 U8473 ( .B1(n14011), .B2(n14047), .A(n14048), .ZN(n14046) );
  AOI211_X1 U8472 ( .C1(n14045), .C2(n14005), .A(n14015), .B(n14046), .ZN(
        n14043) );
  NAND4_X1 U8471 ( .A1(n14041), .A2(n14042), .A3(n14043), .A4(n14021), .ZN(
        \pipeline/cu_pipeline/N103 ) );
  NOR2_X1 U11783 ( .A1(n16993), .A2(n16593), .ZN(\DataMem/N1941 ) );
  NOR2_X1 U11748 ( .A1(n16993), .A2(n16592), .ZN(\DataMem/N2005 ) );
  NOR2_X1 U11889 ( .A1(n16995), .A2(n17651), .ZN(\DataMem/N1745 ) );
  AOI22_X1 U11527 ( .A1(n17660), .A2(\DataMem/Mem[7][23] ), .B1(n17530), .B2(
        \DataMem/Mem[6][23] ), .ZN(n16861) );
  AOI22_X1 U11526 ( .A1(n17531), .A2(\DataMem/Mem[5][23] ), .B1(n16822), .B2(
        \DataMem/Mem[4][23] ), .ZN(n16862) );
  AOI22_X1 U11525 ( .A1(n17122), .A2(\DataMem/Mem[3][23] ), .B1(n16820), .B2(
        \DataMem/Mem[2][23] ), .ZN(n16863) );
  AOI22_X1 U11524 ( .A1(n17124), .A2(\DataMem/Mem[1][23] ), .B1(n17125), .B2(
        \DataMem/Mem[0][23] ), .ZN(n16864) );
  NOR2_X1 U11522 ( .A1(n17155), .A2(n16860), .ZN(\DataMem/N2230 ) );
  NOR2_X1 U11925 ( .A1(n16988), .A2(n16597), .ZN(\DataMem/N1695 ) );
  NOR2_X1 U11804 ( .A1(n16980), .A2(n17655), .ZN(\DataMem/N1903 ) );
  NOR2_X1 U11666 ( .A1(n16980), .A2(n17661), .ZN(\DataMem/N2159 ) );
  NOR2_X1 U11882 ( .A1(n16988), .A2(n16596), .ZN(\DataMem/N1759 ) );
  NOR2_X1 U11939 ( .A1(n16995), .A2(n17650), .ZN(\DataMem/N1681 ) );
  NOR2_X1 U11847 ( .A1(n16988), .A2(n16595), .ZN(\DataMem/N1823 ) );
  NOR2_X1 U11839 ( .A1(n16980), .A2(n17654), .ZN(\DataMem/N1839 ) );
  AOI22_X1 U11479 ( .A1(n17659), .A2(\DataMem/Mem[7][31] ), .B1(n16824), .B2(
        \DataMem/Mem[6][31] ), .ZN(n16813) );
  AOI22_X1 U11478 ( .A1(n16821), .A2(\DataMem/Mem[5][31] ), .B1(n16822), .B2(
        \DataMem/Mem[4][31] ), .ZN(n16814) );
  AOI22_X1 U11477 ( .A1(n17122), .A2(\DataMem/Mem[3][31] ), .B1(n17652), .B2(
        \DataMem/Mem[2][31] ), .ZN(n16815) );
  AOI22_X1 U11476 ( .A1(n16817), .A2(\DataMem/Mem[1][31] ), .B1(n17125), .B2(
        \DataMem/Mem[0][31] ), .ZN(n16816) );
  NOR2_X1 U11474 ( .A1(n12766), .A2(n16812), .ZN(\DataMem/N2254 ) );
  NOR2_X1 U11812 ( .A1(n16988), .A2(n16594), .ZN(\DataMem/N1887 ) );
  AOI22_X1 U11569 ( .A1(n17659), .A2(\DataMem/Mem[7][16] ), .B1(n16824), .B2(
        \DataMem/Mem[6][16] ), .ZN(n16896) );
  AOI22_X1 U11568 ( .A1(n16821), .A2(\DataMem/Mem[5][16] ), .B1(n16822), .B2(
        \DataMem/Mem[4][16] ), .ZN(n16897) );
  AOI22_X1 U11567 ( .A1(n17122), .A2(\DataMem/Mem[3][16] ), .B1(n17653), .B2(
        \DataMem/Mem[2][16] ), .ZN(n16898) );
  AOI22_X1 U11566 ( .A1(n17124), .A2(\DataMem/Mem[1][16] ), .B1(n17125), .B2(
        \DataMem/Mem[0][16] ), .ZN(n16899) );
  NOR2_X1 U11564 ( .A1(n17155), .A2(n16895), .ZN(\DataMem/N2209 ) );
  NOR2_X1 U11778 ( .A1(n16988), .A2(n16593), .ZN(\DataMem/N1951 ) );
  NOR2_X1 U11874 ( .A1(n16980), .A2(n17651), .ZN(\DataMem/N1775 ) );
  NOR2_X1 U11743 ( .A1(n16988), .A2(n16592), .ZN(\DataMem/N2015 ) );
  NOR2_X1 U11708 ( .A1(n16988), .A2(n16591), .ZN(\DataMem/N2079 ) );
  NOR2_X1 U11909 ( .A1(n16980), .A2(n17650), .ZN(\DataMem/N1711 ) );
  NOR2_X1 U11674 ( .A1(n16988), .A2(n16590), .ZN(\DataMem/N2143 ) );
  NOR2_X1 U11680 ( .A1(n16994), .A2(n16590), .ZN(\DataMem/N2131 ) );
  AOI22_X1 U11533 ( .A1(n17660), .A2(\DataMem/Mem[7][22] ), .B1(n17530), .B2(
        \DataMem/Mem[6][22] ), .ZN(n16866) );
  AOI22_X1 U11532 ( .A1(n17531), .A2(\DataMem/Mem[5][22] ), .B1(n16822), .B2(
        \DataMem/Mem[4][22] ), .ZN(n16867) );
  AOI22_X1 U11531 ( .A1(n17122), .A2(\DataMem/Mem[3][22] ), .B1(n16820), .B2(
        \DataMem/Mem[2][22] ), .ZN(n16868) );
  AOI22_X1 U11530 ( .A1(n17124), .A2(\DataMem/Mem[1][22] ), .B1(n17125), .B2(
        \DataMem/Mem[0][22] ), .ZN(n16869) );
  NOR2_X1 U11528 ( .A1(n17155), .A2(n16865), .ZN(\DataMem/N2227 ) );
  AOI22_X1 U11928 ( .A1(\pipeline/Forward_sw1_mux ), .A2(
        \pipeline/data_to_RF_from_WB[22] ), .B1(n13797), .B2(n17380), .ZN(
        n16989) );
  NOR2_X1 U11927 ( .A1(n16989), .A2(n16597), .ZN(\DataMem/N1693 ) );
  NOR2_X1 U11883 ( .A1(n16989), .A2(n16596), .ZN(\DataMem/N1757 ) );
  NOR2_X1 U11848 ( .A1(n16989), .A2(n16595), .ZN(\DataMem/N1821 ) );
  NOR2_X1 U11813 ( .A1(n16989), .A2(n16594), .ZN(\DataMem/N1885 ) );
  NOR2_X1 U11929 ( .A1(n16990), .A2(n16597), .ZN(\DataMem/N1691 ) );
  NOR2_X1 U11779 ( .A1(n16989), .A2(n16593), .ZN(\DataMem/N1949 ) );
  NOR2_X1 U11744 ( .A1(n16989), .A2(n16592), .ZN(\DataMem/N2013 ) );
  NOR2_X1 U11714 ( .A1(n16994), .A2(n16591), .ZN(\DataMem/N2067 ) );
  NOR2_X1 U11709 ( .A1(n16989), .A2(n16591), .ZN(\DataMem/N2077 ) );
  NOR2_X1 U11675 ( .A1(n16989), .A2(n16590), .ZN(\DataMem/N2141 ) );
  NOR2_X1 U11784 ( .A1(n16994), .A2(n16593), .ZN(\DataMem/N1939 ) );
  AOI22_X1 U11539 ( .A1(n17660), .A2(\DataMem/Mem[7][21] ), .B1(n17530), .B2(
        \DataMem/Mem[6][21] ), .ZN(n16871) );
  AOI22_X1 U11538 ( .A1(n16821), .A2(\DataMem/Mem[5][21] ), .B1(n16822), .B2(
        \DataMem/Mem[4][21] ), .ZN(n16872) );
  AOI22_X1 U11537 ( .A1(n17122), .A2(\DataMem/Mem[3][21] ), .B1(n16820), .B2(
        \DataMem/Mem[2][21] ), .ZN(n16873) );
  AOI22_X1 U11536 ( .A1(n17124), .A2(\DataMem/Mem[1][21] ), .B1(n17125), .B2(
        \DataMem/Mem[0][21] ), .ZN(n16874) );
  NOR2_X1 U11534 ( .A1(n17155), .A2(n16870), .ZN(\DataMem/N2224 ) );
  NOR2_X1 U11745 ( .A1(n16990), .A2(n16592), .ZN(\DataMem/N2011 ) );
  NOR2_X1 U11884 ( .A1(n16990), .A2(n16596), .ZN(\DataMem/N1755 ) );
  NOR2_X1 U11749 ( .A1(n16994), .A2(n16592), .ZN(\DataMem/N2003 ) );
  NOR2_X1 U11849 ( .A1(n16990), .A2(n16595), .ZN(\DataMem/N1819 ) );
  NOR2_X1 U11814 ( .A1(n16990), .A2(n16594), .ZN(\DataMem/N1883 ) );
  NOR2_X1 U11780 ( .A1(n16990), .A2(n16593), .ZN(\DataMem/N1947 ) );
  NAND2_X1 U8522 ( .A1(\pipeline/MEM_controls_in_MEM[1] ), .A2(n14105), .ZN(
        n14104) );
  OAI22_X1 U8510 ( .A1(n14103), .A2(n14104), .B1(n14092), .B2(n14105), .ZN(
        n14102) );
  OAI211_X1 U8509 ( .C1(\pipeline/WB_controls_in_MEMWB[1] ), .C2(n14093), .A(
        n14090), .B(n14102), .ZN(\pipeline/cu_hazard/N39 ) );
  NOR2_X1 U8457 ( .A1(\pipeline/inst_IFID_DEC[30] ), .A2(n14011), .ZN(n14008)
         );
  NOR4_X1 U8456 ( .A1(n14007), .A2(n14008), .A3(n14009), .A4(n14010), .ZN(
        n14003) );
  NAND2_X1 U8454 ( .A1(n14005), .A2(n13989), .ZN(n14004) );
  NAND4_X1 U8453 ( .A1(n14002), .A2(n14003), .A3(n17704), .A4(n14004), .ZN(
        \pipeline/cu_pipeline/N109 ) );
  AOI21_X1 U8445 ( .B1(n13980), .B2(n13984), .A(n13281), .ZN(
        \pipeline/cu_pipeline/N113 ) );
  NAND2_X1 U8443 ( .A1(n13982), .A2(n13983), .ZN(\pipeline/cu_pipeline/N112 )
         );
  NOR3_X1 U10220 ( .A1(n17347), .A2(n17313), .A3(n14177), .ZN(n14127) );
  NOR2_X1 U10231 ( .A1(\pipeline/stall ), .A2(n15648), .ZN(n15601) );
  NOR2_X1 U11463 ( .A1(\pipeline/RegDst_to_WB[3] ), .A2(
        \pipeline/RegDst_to_WB[4] ), .ZN(n16584) );
  NOR2_X1 U8654 ( .A1(\pipeline/inst_IFID_DEC[29] ), .A2(n14169), .ZN(n14007)
         );
  NOR4_X1 U8633 ( .A1(n14007), .A2(n14009), .A3(n14183), .A4(n14184), .ZN(
        n13980) );
  NOR3_X1 U8615 ( .A1(\pipeline/inst_IFID_DEC[27] ), .A2(n14176), .A3(n14177), 
        .ZN(\pipeline/cu_pipeline/N89 ) );
  NAND2_X1 U9475 ( .A1(n17703), .A2(\pipeline/WB_controls_in_MEMWB[1] ), .ZN(
        n14129) );
  AOI22_X1 U11950 ( .A1(n17744), .A2(\pipeline/data_to_RF_from_WB[11] ), .B1(
        n13818), .B2(n17743), .ZN(n17000) );
  AOI22_X1 U11952 ( .A1(\pipeline/Forward_sw1_mux ), .A2(
        \pipeline/data_to_RF_from_WB[10] ), .B1(n13816), .B2(n17743), .ZN(
        n17001) );
  AOI22_X1 U11948 ( .A1(\pipeline/Forward_sw1_mux ), .A2(
        \pipeline/data_to_RF_from_WB[12] ), .B1(n13812), .B2(n17380), .ZN(
        n16999) );
  AOI22_X1 U11968 ( .A1(n17744), .A2(\pipeline/data_to_RF_from_WB[2] ), .B1(
        n13808), .B2(n17743), .ZN(n17009) );
  AOI22_X1 U11966 ( .A1(n17744), .A2(\pipeline/data_to_RF_from_WB[3] ), .B1(
        n13807), .B2(n17743), .ZN(n17008) );
  AOI22_X1 U11970 ( .A1(\pipeline/Forward_sw1_mux ), .A2(
        \pipeline/data_to_RF_from_WB[1] ), .B1(n13805), .B2(n17743), .ZN(
        n17010) );
  AOI22_X1 U11958 ( .A1(n17744), .A2(\pipeline/data_to_RF_from_WB[7] ), .B1(
        n13830), .B2(n17743), .ZN(n17004) );
  AOI22_X1 U11964 ( .A1(n17744), .A2(\pipeline/data_to_RF_from_WB[4] ), .B1(
        n13835), .B2(n17743), .ZN(n17007) );
  AOI22_X1 U11960 ( .A1(n17744), .A2(\pipeline/data_to_RF_from_WB[6] ), .B1(
        n13828), .B2(n17743), .ZN(n17005) );
  AOI22_X1 U11962 ( .A1(n17744), .A2(\pipeline/data_to_RF_from_WB[5] ), .B1(
        n13831), .B2(n17743), .ZN(n17006) );
  AOI22_X1 U11954 ( .A1(\pipeline/Forward_sw1_mux ), .A2(
        \pipeline/data_to_RF_from_WB[9] ), .B1(n13819), .B2(n17743), .ZN(
        n17002) );
  AOI22_X1 U11912 ( .A1(n17744), .A2(\pipeline/data_to_RF_from_WB[30] ), .B1(
        n13791), .B2(n17380), .ZN(n16981) );
  AOI22_X1 U11956 ( .A1(n17744), .A2(\pipeline/data_to_RF_from_WB[8] ), .B1(
        n13785), .B2(n17743), .ZN(n17003) );
  AOI22_X1 U11914 ( .A1(\pipeline/Forward_sw1_mux ), .A2(
        \pipeline/data_to_RF_from_WB[29] ), .B1(n13792), .B2(n17743), .ZN(
        n16982) );
  AOI22_X1 U11976 ( .A1(n17744), .A2(\pipeline/data_to_RF_from_WB[0] ), .B1(
        n13784), .B2(n17743), .ZN(n17011) );
  AOI22_X1 U11922 ( .A1(n17744), .A2(\pipeline/data_to_RF_from_WB[25] ), .B1(
        n13795), .B2(n17743), .ZN(n16986) );
  AOI22_X1 U11916 ( .A1(n17744), .A2(\pipeline/data_to_RF_from_WB[28] ), .B1(
        n13787), .B2(n17380), .ZN(n16983) );
  AOI22_X1 U11924 ( .A1(n17744), .A2(\pipeline/data_to_RF_from_WB[24] ), .B1(
        n13786), .B2(n17743), .ZN(n16987) );
  AOI22_X1 U11944 ( .A1(n17744), .A2(\pipeline/data_to_RF_from_WB[14] ), .B1(
        n13788), .B2(n17380), .ZN(n16997) );
  AOI22_X1 U11942 ( .A1(\pipeline/Forward_sw1_mux ), .A2(
        \pipeline/data_to_RF_from_WB[15] ), .B1(n13789), .B2(n17380), .ZN(
        n16996) );
  AOI22_X1 U11930 ( .A1(n17744), .A2(\pipeline/data_to_RF_from_WB[21] ), .B1(
        n13798), .B2(n17380), .ZN(n16990) );
  AOI22_X1 U11938 ( .A1(\pipeline/Forward_sw1_mux ), .A2(
        \pipeline/data_to_RF_from_WB[17] ), .B1(n13802), .B2(n17380), .ZN(
        n16994) );
  AOI22_X1 U11932 ( .A1(n17744), .A2(\pipeline/data_to_RF_from_WB[20] ), .B1(
        n13799), .B2(n17380), .ZN(n16991) );
  AOI22_X1 U11926 ( .A1(n17744), .A2(\pipeline/data_to_RF_from_WB[23] ), .B1(
        n13796), .B2(n17743), .ZN(n16988) );
  NAND3_X1 U12241 ( .A1(\pipeline/RegDst_to_WB[3] ), .A2(
        \pipeline/RegDst_to_WB[4] ), .A3(n17643), .ZN(n16589) );
  NAND3_X1 U12234 ( .A1(\pipeline/RegDst_to_WB[4] ), .A2(n17643), .A3(n17385), 
        .ZN(n16588) );
  NAND3_X1 U12233 ( .A1(\pipeline/RegDst_to_WB[3] ), .A2(n17643), .A3(n17386), 
        .ZN(n16587) );
  NOR2_X1 U10247 ( .A1(\pipeline/inst_IFID_DEC[31] ), .A2(n17348), .ZN(n14049)
         );
  NOR2_X1 U10244 ( .A1(n14186), .A2(n14059), .ZN(n14126) );
  NOR2_X1 U10240 ( .A1(\pipeline/inst_IFID_DEC[30] ), .A2(
        \pipeline/inst_IFID_DEC[26] ), .ZN(n13993) );
  NOR2_X1 U9893 ( .A1(n13281), .A2(\pipeline/EXE_controls_in_EXEcute [5]), 
        .ZN(n14995) );
  NAND2_X1 U9871 ( .A1(\pipeline/EXE_controls_in_EXEcute [2]), .A2(n15573), 
        .ZN(n14981) );
  NAND2_X1 U9389 ( .A1(\pipeline/stageD/offset_jump_sign_ext [18]), .A2(
        \pipeline/stageD/offset_jump_sign_ext [17]), .ZN(n14863) );
  NAND2_X1 U9383 ( .A1(\pipeline/stageD/offset_jump_sign_ext [18]), .A2(n17329), .ZN(n14865) );
  NAND2_X1 U9371 ( .A1(\pipeline/stageD/offset_jump_sign_ext [17]), .A2(n17408), .ZN(n14864) );
  NOR2_X1 U11426 ( .A1(n16785), .A2(n16786), .ZN(n16778) );
  NOR2_X1 U10212 ( .A1(n15827), .A2(n15828), .ZN(n15606) );
  NAND3_X1 U11978 ( .A1(\pipeline/stageD/offset_to_jump_temp [15]), .A2(
        \pipeline/EXE_controls_in_IDEX[8] ), .A3(n13967), .ZN(n13969) );
  OAI21_X1 U8431 ( .B1(n13967), .B2(n17328), .A(n13969), .ZN(
        \pipeline/stageD/offset_to_jump_temp [30]) );
  NAND2_X1 U10922 ( .A1(\pipeline/WB_controls_in_MEMWB[1] ), .A2(n14103), .ZN(
        n15827) );
  OAI21_X1 U10237 ( .B1(n15839), .B2(n15840), .A(n15841), .ZN(n15838) );
  NOR2_X1 U10213 ( .A1(n15829), .A2(n15828), .ZN(n15605) );
  NOR2_X1 U10902 ( .A1(n16546), .A2(n16532), .ZN(n15930) );
  NOR2_X1 U10901 ( .A1(n16545), .A2(n16532), .ZN(n15931) );
  NOR2_X1 U10899 ( .A1(n16530), .A2(n16540), .ZN(n15928) );
  NOR2_X1 U10898 ( .A1(n16530), .A2(n16539), .ZN(n15929) );
  NOR2_X1 U10896 ( .A1(n16529), .A2(n16540), .ZN(n15926) );
  NOR2_X1 U10895 ( .A1(n16529), .A2(n16539), .ZN(n15927) );
  NOR2_X1 U10893 ( .A1(n16532), .A2(n16540), .ZN(n15924) );
  NOR2_X1 U10892 ( .A1(n16532), .A2(n16539), .ZN(n15925) );
  NOR4_X1 U10929 ( .A1(n16560), .A2(n16561), .A3(n16562), .A4(n16563), .ZN(
        n15830) );
  NOR2_X1 U10915 ( .A1(n16546), .A2(n16530), .ZN(n15940) );
  NOR2_X1 U10914 ( .A1(n16530), .A2(n16545), .ZN(n15941) );
  NAND2_X1 U10912 ( .A1(\pipeline/stageD/offset_jump_sign_ext [23]), .A2(
        n17317), .ZN(n16529) );
  NOR2_X1 U10911 ( .A1(n16546), .A2(n16529), .ZN(n15938) );
  NOR2_X1 U10910 ( .A1(n16545), .A2(n16529), .ZN(n15939) );
  NOR2_X1 U10889 ( .A1(n16527), .A2(n16540), .ZN(n15918) );
  NOR2_X1 U10885 ( .A1(n16532), .A2(n16531), .ZN(n15917) );
  NOR2_X1 U10883 ( .A1(n16533), .A2(n16529), .ZN(n15914) );
  NOR2_X1 U10880 ( .A1(n16533), .A2(n16530), .ZN(n15912) );
  OAI21_X1 U10249 ( .B1(n15830), .B2(n15842), .A(n15843), .ZN(n15839) );
  NAND2_X1 U10916 ( .A1(\pipeline/stageD/offset_jump_sign_ext [22]), .A2(
        \pipeline/stageD/offset_jump_sign_ext [23]), .ZN(n16530) );
  NAND2_X1 U10908 ( .A1(n17317), .A2(n17383), .ZN(n16527) );
  NOR2_X1 U10907 ( .A1(n16527), .A2(n16533), .ZN(n15935) );
  NOR2_X1 U10906 ( .A1(n16527), .A2(n16546), .ZN(n15936) );
  NOR2_X1 U10905 ( .A1(n16527), .A2(n16545), .ZN(n15937) );
  NAND2_X1 U10903 ( .A1(\pipeline/stageD/offset_jump_sign_ext [22]), .A2(
        n17383), .ZN(n16532) );
  NOR2_X1 U10876 ( .A1(n16529), .A2(n16534), .ZN(n15906) );
  NOR2_X1 U10872 ( .A1(n16532), .A2(n16528), .ZN(n15905) );
  NOR2_X1 U10869 ( .A1(n16530), .A2(n16528), .ZN(n15903) );
  OAI21_X1 U10233 ( .B1(n15834), .B2(n14947), .A(n17703), .ZN(n15648) );
  AOI21_X1 U10236 ( .B1(n13979), .B2(n15646), .A(n15838), .ZN(n15834) );
  INV_X1 U8441 ( .A(n13979), .ZN(n13967) );
  INV_X1 U10936 ( .A(n16555), .ZN(n16560) );
  INV_X1 U10766 ( .A(n15827), .ZN(n15832) );
  INV_X1 U10746 ( .A(n14945), .ZN(n15772) );
  INV_X1 U10726 ( .A(n14883), .ZN(n15688) );
  INV_X1 U10260 ( .A(n15886), .ZN(n15842) );
  INV_X1 U10239 ( .A(n13993), .ZN(n14176) );
  INV_X1 U10224 ( .A(n15834), .ZN(n15833) );
  NAND2_X1 U10218 ( .A1(n15833), .A2(n14127), .ZN(n15828) );
  INV_X1 U10214 ( .A(n15830), .ZN(n15829) );
  INV_X1 U11317 ( .A(n15427), .ZN(n15426) );
  OAI21_X1 U11313 ( .B1(n17662), .B2(n17344), .A(n16729), .ZN(
        \pipeline/stageE/input1_to_ALU [13]) );
  INV_X1 U11218 ( .A(\pipeline/stageE/input1_to_ALU [4]), .ZN(n15564) );
  OR2_X1 U11217 ( .A1(n16683), .A2(n15564), .ZN(n15569) );
  INV_X1 U11209 ( .A(n15538), .ZN(n15537) );
  OR2_X1 U11201 ( .A1(\pipeline/stageE/input1_to_ALU [6]), .A2(n16676), .ZN(
        n15527) );
  INV_X1 U11289 ( .A(n15498), .ZN(n15505) );
  OR2_X1 U11287 ( .A1(\pipeline/stageE/input1_to_ALU [8]), .A2(n16672), .ZN(
        n15509) );
  INV_X1 U11187 ( .A(n15492), .ZN(n15491) );
  INV_X1 U11184 ( .A(n15477), .ZN(n15495) );
  INV_X1 U11174 ( .A(n15435), .ZN(n15442) );
  INV_X1 U11167 ( .A(n15431), .ZN(n15446) );
  INV_X1 U11164 ( .A(n15414), .ZN(n15432) );
  INV_X1 U11158 ( .A(n15411), .ZN(n15410) );
  INV_X1 U11151 ( .A(n15400), .ZN(n15413) );
  INV_X1 U11134 ( .A(n15363), .ZN(n15362) );
  INV_X1 U11131 ( .A(n16632), .ZN(n15367) );
  INV_X1 U11123 ( .A(n15372), .ZN(n15379) );
  OR2_X1 U11121 ( .A1(\pipeline/stageE/EXE_ALU/alu_shift/C48/A[16] ), .A2(
        n15369), .ZN(n15383) );
  INV_X1 U11111 ( .A(n15331), .ZN(n15330) );
  OAI21_X1 U11335 ( .B1(n17105), .B2(n17322), .A(n16738), .ZN(
        \pipeline/stageE/input1_to_ALU [20]) );
  INV_X1 U11353 ( .A(n15279), .ZN(n15278) );
  OAI21_X1 U11089 ( .B1(n17662), .B2(n17324), .A(n16618), .ZN(
        \pipeline/stageE/input1_to_ALU [24]) );
  INV_X1 U11083 ( .A(n15246), .ZN(n15245) );
  INV_X1 U11081 ( .A(n15249), .ZN(n16613) );
  OAI21_X1 U11368 ( .B1(n17662), .B2(n17427), .A(n16754), .ZN(
        \pipeline/stageE/input1_to_ALU [25]) );
  OR2_X1 U11390 ( .A1(n16611), .A2(\pipeline/stageE/input1_to_ALU [28]), .ZN(
        n15166) );
  INV_X1 U9653 ( .A(n15221), .ZN(n15219) );
  INV_X1 U9703 ( .A(n15301), .ZN(n15300) );
  INV_X1 U9806 ( .A(n15476), .ZN(n15462) );
  INV_X1 U9859 ( .A(n15540), .ZN(n15555) );
  INV_X1 U9897 ( .A(n15056), .ZN(n15594) );
  INV_X1 U9511 ( .A(n15055), .ZN(n15054) );
  INV_X1 U9717 ( .A(n15297), .ZN(n15320) );
  INV_X1 U11403 ( .A(n15169), .ZN(n15176) );
  INV_X1 U9611 ( .A(n15162), .ZN(n15145) );
  INV_X1 U11411 ( .A(n15150), .ZN(n15157) );
  INV_X1 U11063 ( .A(n15134), .ZN(n15133) );
  INV_X1 U10052 ( .A(n14889), .ZN(n15692) );
  INV_X1 U10058 ( .A(n14891), .ZN(n15697) );
  INV_X1 U9889 ( .A(n15588), .ZN(n15573) );
  INV_X1 U9867 ( .A(n14949), .ZN(n14993) );
  INV_X1 U10064 ( .A(n14893), .ZN(n15702) );
  INV_X1 U9630 ( .A(n15182), .ZN(n15189) );
  INV_X1 U10070 ( .A(n14895), .ZN(n15707) );
  INV_X1 U9640 ( .A(n15202), .ZN(n15201) );
  INV_X1 U9650 ( .A(n15216), .ZN(n15215) );
  INV_X1 U10076 ( .A(n14897), .ZN(n15712) );
  INV_X1 U9677 ( .A(n15261), .ZN(n15260) );
  INV_X1 U9659 ( .A(n15224), .ZN(n15231) );
  INV_X1 U10082 ( .A(n14899), .ZN(n15717) );
  INV_X1 U9711 ( .A(n15312), .ZN(n15311) );
  INV_X1 U9699 ( .A(n15285), .ZN(n15292) );
  INV_X1 U9792 ( .A(n15449), .ZN(n15456) );
  INV_X1 U9732 ( .A(n15346), .ZN(n15345) );
  INV_X1 U9776 ( .A(\pipeline/stageE/input1_to_ALU [13]), .ZN(n15425) );
  INV_X1 U9759 ( .A(n15386), .ZN(n15393) );
  INV_X1 U10088 ( .A(n14901), .ZN(n15722) );
  INV_X1 U9856 ( .A(n15553), .ZN(n15552) );
  INV_X1 U9805 ( .A(n15474), .ZN(n15473) );
  INV_X1 U9832 ( .A(n15512), .ZN(n15519) );
  INV_X1 U10094 ( .A(n14903), .ZN(n15727) );
  INV_X1 U9980 ( .A(n15653), .ZN(n3957) );
  INV_X1 U9972 ( .A(n15649), .ZN(n3961) );
  INV_X1 U9968 ( .A(n15645), .ZN(n3963) );
  INV_X1 U9960 ( .A(n15641), .ZN(n3967) );
  INV_X1 U9976 ( .A(n15651), .ZN(n3959) );
  INV_X1 U9962 ( .A(n15642), .ZN(n3966) );
  INV_X1 U10144 ( .A(n15768), .ZN(n3881) );
  INV_X1 U10155 ( .A(n15778), .ZN(n3877) );
  INV_X1 U10066 ( .A(n15703), .ZN(n3907) );
  INV_X1 U9940 ( .A(n15631), .ZN(n3977) );
  INV_X1 U9964 ( .A(n15643), .ZN(n3965) );
  INV_X1 U10054 ( .A(n15693), .ZN(n3911) );
  INV_X1 U10197 ( .A(n15813), .ZN(n3863) );
  INV_X1 U10173 ( .A(n15793), .ZN(n3871) );
  INV_X1 U9930 ( .A(n15626), .ZN(n3982) );
  INV_X1 U10090 ( .A(n15723), .ZN(n3899) );
  INV_X1 U10108 ( .A(n15738), .ZN(n3893) );
  INV_X1 U9952 ( .A(n15637), .ZN(n3971) );
  INV_X1 U10167 ( .A(n15788), .ZN(n3873) );
  INV_X1 U9928 ( .A(n15625), .ZN(n3983) );
  INV_X1 U10078 ( .A(n15713), .ZN(n3903) );
  INV_X1 U10138 ( .A(n15763), .ZN(n3883) );
  INV_X1 U9904 ( .A(n15599), .ZN(n3992) );
  INV_X1 U9950 ( .A(n15636), .ZN(n3972) );
  INV_X1 U10161 ( .A(n15783), .ZN(n3875) );
  INV_X1 U10229 ( .A(n15837), .ZN(n3855) );
  INV_X1 U9956 ( .A(n15639), .ZN(n3969) );
  INV_X1 U10209 ( .A(n15823), .ZN(n3859) );
  INV_X1 U9958 ( .A(n15640), .ZN(n3968) );
  INV_X1 U10126 ( .A(n15753), .ZN(n3887) );
  INV_X1 U10120 ( .A(n15748), .ZN(n3889) );
  INV_X1 U10102 ( .A(n15733), .ZN(n3895) );
  INV_X1 U9938 ( .A(n15630), .ZN(n3978) );
  INV_X1 U9946 ( .A(n15634), .ZN(n3974) );
  INV_X1 U9942 ( .A(n15632), .ZN(n3976) );
  INV_X1 U10072 ( .A(n15708), .ZN(n3905) );
  INV_X1 U10096 ( .A(n15728), .ZN(n3897) );
  INV_X1 U9922 ( .A(n15622), .ZN(n3986) );
  INV_X1 U9932 ( .A(n15627), .ZN(n3981) );
  INV_X1 U9944 ( .A(n15633), .ZN(n3975) );
  INV_X1 U10060 ( .A(n15698), .ZN(n3909) );
  INV_X1 U10203 ( .A(n15818), .ZN(n3861) );
  INV_X1 U10191 ( .A(n15808), .ZN(n3865) );
  INV_X1 U10185 ( .A(n15803), .ZN(n3867) );
  INV_X1 U10225 ( .A(n15835), .ZN(n3857) );
  INV_X1 U10149 ( .A(n15773), .ZN(n3879) );
  INV_X1 U9924 ( .A(n15623), .ZN(n3985) );
  INV_X1 U9954 ( .A(n15638), .ZN(n3970) );
  INV_X1 U9948 ( .A(n15635), .ZN(n3973) );
  INV_X1 U10100 ( .A(n14905), .ZN(n15732) );
  AND2_X1 U10049 ( .A1(n15600), .A2(n13937), .ZN(n3923) );
  INV_X1 U10201 ( .A(n14921), .ZN(n15817) );
  INV_X1 U10142 ( .A(n14929), .ZN(n15767) );
  INV_X1 U10112 ( .A(n14909), .ZN(n15742) );
  INV_X1 U10124 ( .A(n14915), .ZN(n15752) );
  INV_X1 U10153 ( .A(n14939), .ZN(n15777) );
  INV_X1 U9908 ( .A(n14913), .ZN(n15609) );
  INV_X1 U10195 ( .A(n14925), .ZN(n15812) );
  INV_X1 U10165 ( .A(n14937), .ZN(n15787) );
  INV_X1 U10207 ( .A(n14941), .ZN(n15822) );
  INV_X1 U10132 ( .A(n15758), .ZN(n3885) );
  INV_X1 U10114 ( .A(n15743), .ZN(n3891) );
  INV_X1 U9936 ( .A(n15629), .ZN(n3979) );
  INV_X1 U10227 ( .A(n15836), .ZN(n3856) );
  INV_X1 U10177 ( .A(n14933), .ZN(n15797) );
  INV_X1 U10136 ( .A(n14919), .ZN(n15762) );
  INV_X1 U10106 ( .A(n14907), .ZN(n15737) );
  INV_X1 U10171 ( .A(n14935), .ZN(n15792) );
  INV_X1 U10159 ( .A(n14931), .ZN(n15782) );
  INV_X1 U10118 ( .A(n14911), .ZN(n15747) );
  INV_X1 U10216 ( .A(n14943), .ZN(n15831) );
  INV_X1 U10183 ( .A(n14923), .ZN(n15802) );
  INV_X1 U10130 ( .A(n14917), .ZN(n15757) );
  INV_X1 U10189 ( .A(n14927), .ZN(n15807) );
  INV_X1 U9966 ( .A(n15644), .ZN(n3964) );
  INV_X1 U9934 ( .A(n15628), .ZN(n3980) );
  INV_X1 U9926 ( .A(n15624), .ZN(n3984) );
  INV_X1 U9910 ( .A(n15612), .ZN(n3990) );
  INV_X1 U10179 ( .A(n15798), .ZN(n3869) );
  INV_X1 U10084 ( .A(n15718), .ZN(n3901) );
  INV_X1 U9456 ( .A(n14947), .ZN(n14025) );
  INV_X1 U8652 ( .A(n13998), .ZN(n14001) );
  INV_X1 U8646 ( .A(n14011), .ZN(n14185) );
  AND2_X1 U8623 ( .A1(n17412), .A2(n14179), .ZN(n14044) );
  INV_X1 U8593 ( .A(n14165), .ZN(\pipeline/MEMWB_Stage/N12 ) );
  INV_X1 U8595 ( .A(n14166), .ZN(\pipeline/MEMWB_Stage/N11 ) );
  INV_X1 U8565 ( .A(n14151), .ZN(\pipeline/MEMWB_Stage/N26 ) );
  INV_X1 U8569 ( .A(n14153), .ZN(\pipeline/MEMWB_Stage/N24 ) );
  INV_X1 U8547 ( .A(n14142), .ZN(\pipeline/MEMWB_Stage/N35 ) );
  INV_X1 U8583 ( .A(n14160), .ZN(\pipeline/MEMWB_Stage/N17 ) );
  INV_X1 U8539 ( .A(n14138), .ZN(\pipeline/MEMWB_Stage/N39 ) );
  INV_X1 U8571 ( .A(n14154), .ZN(\pipeline/MEMWB_Stage/N23 ) );
  INV_X1 U8533 ( .A(n14133), .ZN(\pipeline/MEMWB_Stage/N42 ) );
  INV_X1 U8545 ( .A(n14141), .ZN(\pipeline/MEMWB_Stage/N36 ) );
  INV_X1 U8549 ( .A(n14143), .ZN(\pipeline/MEMWB_Stage/N34 ) );
  INV_X1 U8587 ( .A(n14162), .ZN(\pipeline/MEMWB_Stage/N15 ) );
  INV_X1 U8589 ( .A(n14163), .ZN(\pipeline/MEMWB_Stage/N14 ) );
  INV_X1 U8579 ( .A(n14158), .ZN(\pipeline/MEMWB_Stage/N19 ) );
  INV_X1 U8581 ( .A(n14159), .ZN(\pipeline/MEMWB_Stage/N18 ) );
  INV_X1 U8551 ( .A(n14144), .ZN(\pipeline/MEMWB_Stage/N33 ) );
  INV_X1 U8591 ( .A(n14164), .ZN(\pipeline/MEMWB_Stage/N13 ) );
  INV_X1 U8577 ( .A(n14157), .ZN(\pipeline/MEMWB_Stage/N20 ) );
  INV_X1 U8553 ( .A(n14145), .ZN(\pipeline/MEMWB_Stage/N32 ) );
  INV_X1 U8573 ( .A(n14155), .ZN(\pipeline/MEMWB_Stage/N22 ) );
  INV_X1 U8559 ( .A(n14148), .ZN(\pipeline/MEMWB_Stage/N29 ) );
  INV_X1 U8555 ( .A(n14146), .ZN(\pipeline/MEMWB_Stage/N31 ) );
  INV_X1 U8535 ( .A(n14136), .ZN(\pipeline/MEMWB_Stage/N41 ) );
  INV_X1 U8537 ( .A(n14137), .ZN(\pipeline/MEMWB_Stage/N40 ) );
  INV_X1 U8541 ( .A(n14139), .ZN(\pipeline/MEMWB_Stage/N38 ) );
  INV_X1 U8557 ( .A(n14147), .ZN(\pipeline/MEMWB_Stage/N30 ) );
  INV_X1 U8543 ( .A(n14140), .ZN(\pipeline/MEMWB_Stage/N37 ) );
  INV_X1 U8567 ( .A(n14152), .ZN(\pipeline/MEMWB_Stage/N25 ) );
  INV_X1 U8585 ( .A(n14161), .ZN(\pipeline/MEMWB_Stage/N16 ) );
  INV_X1 U8561 ( .A(n14149), .ZN(\pipeline/MEMWB_Stage/N28 ) );
  INV_X1 U8563 ( .A(n14150), .ZN(\pipeline/MEMWB_Stage/N27 ) );
  INV_X1 U8575 ( .A(n14156), .ZN(\pipeline/MEMWB_Stage/N21 ) );
  AND2_X1 U8604 ( .A1(n14167), .A2(\pipeline/EXE_controls_in_IDEX[2] ), .ZN(
        \pipeline/IDEX_Stage/N95 ) );
  AND2_X1 U8601 ( .A1(n14167), .A2(\pipeline/EXE_controls_in_IDEX[5] ), .ZN(
        \pipeline/IDEX_Stage/N98 ) );
  AND2_X1 U8602 ( .A1(n14167), .A2(\pipeline/EXE_controls_in_IDEX[4] ), .ZN(
        \pipeline/IDEX_Stage/N97 ) );
  AND2_X1 U9458 ( .A1(n14167), .A2(\pipeline/EXE_controls_in_IDEX[7] ), .ZN(
        \pipeline/IDEX_Stage/N100 ) );
  AND2_X1 U9457 ( .A1(n14167), .A2(\pipeline/EXE_controls_in_IDEX[8] ), .ZN(
        \pipeline/IDEX_Stage/N101 ) );
  AND2_X1 U8600 ( .A1(n14167), .A2(\pipeline/EXE_controls_in_IDEX[6] ), .ZN(
        \pipeline/IDEX_Stage/N99 ) );
  AND2_X1 U8603 ( .A1(n14167), .A2(\pipeline/EXE_controls_in_IDEX[3] ), .ZN(
        \pipeline/IDEX_Stage/N96 ) );
  AND2_X1 U8656 ( .A1(n14167), .A2(\pipeline/WB_controls_in_IDEX[0] ), .ZN(
        \pipeline/IDEX_Stage/N89 ) );
  AND2_X1 U8605 ( .A1(n14167), .A2(\pipeline/EXE_controls_in_IDEX[1] ), .ZN(
        \pipeline/IDEX_Stage/N94 ) );
  AND2_X1 U8606 ( .A1(n14167), .A2(\pipeline/EXE_controls_in_IDEX[0] ), .ZN(
        \pipeline/IDEX_Stage/N93 ) );
  INV_X1 U8610 ( .A(n14123), .ZN(n13981) );
  INV_X1 U8599 ( .A(n14129), .ZN(\pipeline/MEMWB_Stage/N10 ) );
  AND2_X1 U8532 ( .A1(\pipeline/regDst_to_mem[0] ), .A2(
        \pipeline/MEMWB_Stage/N10 ), .ZN(\pipeline/MEMWB_Stage/N43 ) );
  INV_X1 U9477 ( .A(n14120), .ZN(n14101) );
  AND2_X1 U9682 ( .A1(n13936), .A2(n17705), .ZN(\pipeline/EXMEM_stage/N3 ) );
  AND2_X1 U9542 ( .A1(\pipeline/MEM_controls_in_EXMEM[1] ), .A2(n17705), .ZN(
        \pipeline/EXMEM_stage/N6 ) );
  NOR3_X2 U11975 ( .A1(addr_to_dataRam[4]), .A2(addr_to_dataRam[2]), .A3(
        addr_to_dataRam[3]), .ZN(n16818) );
  NOR3_X2 U11907 ( .A1(addr_to_dataRam[4]), .A2(addr_to_dataRam[3]), .A3(
        n17012), .ZN(n16817) );
  AND4_X1 U11595 ( .A1(n16921), .A2(n16922), .A3(n16923), .A4(n16924), .ZN(
        n16920) );
  AND4_X1 U11589 ( .A1(n16916), .A2(n16917), .A3(n16918), .A4(n16919), .ZN(
        n16915) );
  AND4_X1 U11649 ( .A1(n16966), .A2(n16967), .A3(n16968), .A4(n16969), .ZN(
        n16965) );
  AND4_X1 U11643 ( .A1(n16961), .A2(n16962), .A3(n16963), .A4(n16964), .ZN(
        n16960) );
  AND4_X1 U11637 ( .A1(n16956), .A2(n16957), .A3(n16958), .A4(n16959), .ZN(
        n16955) );
  AND4_X1 U11601 ( .A1(n16926), .A2(n16927), .A3(n16928), .A4(n16929), .ZN(
        n16925) );
  AND4_X1 U11619 ( .A1(n16941), .A2(n16942), .A3(n16943), .A4(n16944), .ZN(
        n16940) );
  AND4_X1 U11631 ( .A1(n16951), .A2(n16952), .A3(n16953), .A4(n16954), .ZN(
        n16950) );
  AND4_X1 U11607 ( .A1(n16931), .A2(n16932), .A3(n16933), .A4(n16934), .ZN(
        n16930) );
  AND4_X1 U11655 ( .A1(n16971), .A2(n16972), .A3(n16973), .A4(n16974), .ZN(
        n16970) );
  AND4_X1 U11625 ( .A1(n16946), .A2(n16947), .A3(n16948), .A4(n16949), .ZN(
        n16945) );
  AND4_X1 U11487 ( .A1(n16831), .A2(n16832), .A3(n16833), .A4(n16834), .ZN(
        n16830) );
  AND4_X1 U11613 ( .A1(n16936), .A2(n16937), .A3(n16938), .A4(n16939), .ZN(
        n16935) );
  AND4_X1 U11499 ( .A1(n16841), .A2(n16842), .A3(n16843), .A4(n16844), .ZN(
        n16840) );
  AND4_X1 U11505 ( .A1(n16846), .A2(n16847), .A3(n16848), .A4(n16849), .ZN(
        n16845) );
  AND4_X1 U11661 ( .A1(n16976), .A2(n16977), .A3(n16978), .A4(n16979), .ZN(
        n16975) );
  AND4_X1 U11511 ( .A1(n16851), .A2(n16852), .A3(n16853), .A4(n16854), .ZN(
        n16850) );
  AND4_X1 U11577 ( .A1(n16906), .A2(n16907), .A3(n16908), .A4(n16909), .ZN(
        n16905) );
  AND4_X1 U11571 ( .A1(n16901), .A2(n16902), .A3(n16903), .A4(n16904), .ZN(
        n16900) );
  AND4_X1 U11517 ( .A1(n16856), .A2(n16857), .A3(n16858), .A4(n16859), .ZN(
        n16855) );
  AND4_X1 U11583 ( .A1(n16911), .A2(n16912), .A3(n16913), .A4(n16914), .ZN(
        n16910) );
  AND4_X1 U11481 ( .A1(n16826), .A2(n16827), .A3(n16828), .A4(n16829), .ZN(
        n16825) );
  AND4_X1 U11493 ( .A1(n16836), .A2(n16837), .A3(n16838), .A4(n16839), .ZN(
        n16835) );
  AND4_X1 U11541 ( .A1(n16876), .A2(n16877), .A3(n16878), .A4(n16879), .ZN(
        n16875) );
  AND4_X1 U11547 ( .A1(n16881), .A2(n16882), .A3(n16883), .A4(n16884), .ZN(
        n16880) );
  AND4_X1 U11559 ( .A1(n16891), .A2(n16892), .A3(n16893), .A4(n16894), .ZN(
        n16890) );
  INV_X1 U8525 ( .A(n14094), .ZN(n14091) );
  AND3_X1 U8485 ( .A1(n14005), .A2(n14067), .A3(n17350), .ZN(n14033) );
  AND2_X1 U8466 ( .A1(n13981), .A2(n14030), .ZN(n14002) );
  AND2_X1 U8474 ( .A1(n14051), .A2(n14033), .ZN(n14015) );
  INV_X1 U8455 ( .A(n14006), .ZN(n13989) );
  INV_X1 U8496 ( .A(\pipeline/cu_pipeline/N89 ), .ZN(n13984) );
  AND4_X1 U11553 ( .A1(n16886), .A2(n16887), .A3(n16888), .A4(n16889), .ZN(
        n16885) );
  INV_X1 U8489 ( .A(n14005), .ZN(n14012) );
  INV_X1 U8480 ( .A(n14061), .ZN(n14020) );
  INV_X1 U8458 ( .A(n13988), .ZN(\pipeline/cu_pipeline/N108 ) );
  INV_X1 U8462 ( .A(n14022), .ZN(n14018) );
  INV_X1 U8470 ( .A(n14040), .ZN(n14034) );
  AND4_X1 U11523 ( .A1(n16861), .A2(n16862), .A3(n16863), .A4(n16864), .ZN(
        n16860) );
  AND4_X1 U11475 ( .A1(n16813), .A2(n16814), .A3(n16815), .A4(n16816), .ZN(
        n16812) );
  AND4_X1 U11565 ( .A1(n16896), .A2(n16897), .A3(n16898), .A4(n16899), .ZN(
        n16895) );
  AND4_X1 U11529 ( .A1(n16866), .A2(n16867), .A3(n16868), .A4(n16869), .ZN(
        n16865) );
  AND4_X1 U11535 ( .A1(n16871), .A2(n16872), .A3(n16873), .A4(n16874), .ZN(
        n16870) );
  INV_X1 U8523 ( .A(n14093), .ZN(n14105) );
  INV_X1 U8444 ( .A(\pipeline/cu_pipeline/N113 ), .ZN(n13982) );
  DFF_X2 \pipeline/IFID_stage/Instr_out_IFID_reg[0]  ( .D(n3987), .CK(Clk), 
        .Q(net175543), .QN(n17076) );
  INV_X1 \pipeline/stageF/PC_plus4/add_26/U56  ( .A(addr_to_iram[2]), .ZN(
        \pipeline/stageF/PC_plus4/N9 ) );
  AND2_X1 \pipeline/stageF/PC_plus4/add_26/U54  ( .A1(
        \pipeline/stageF/PC_plus4/add_26/carry[28] ), .A2(addr_to_iram[28]), 
        .ZN(\pipeline/stageF/PC_plus4/add_26/carry[29] ) );
  AND2_X1 \pipeline/stageF/PC_plus4/add_26/U52  ( .A1(
        \pipeline/stageF/PC_plus4/add_26/carry[27] ), .A2(addr_to_iram[27]), 
        .ZN(\pipeline/stageF/PC_plus4/add_26/carry[28] ) );
  AND2_X1 \pipeline/stageF/PC_plus4/add_26/U50  ( .A1(
        \pipeline/stageF/PC_plus4/add_26/carry[26] ), .A2(addr_to_iram[26]), 
        .ZN(\pipeline/stageF/PC_plus4/add_26/carry[27] ) );
  AND2_X1 \pipeline/stageF/PC_plus4/add_26/U48  ( .A1(
        \pipeline/stageF/PC_plus4/add_26/carry[25] ), .A2(addr_to_iram[25]), 
        .ZN(\pipeline/stageF/PC_plus4/add_26/carry[26] ) );
  AND2_X1 \pipeline/stageF/PC_plus4/add_26/U46  ( .A1(
        \pipeline/stageF/PC_plus4/add_26/carry[24] ), .A2(addr_to_iram[24]), 
        .ZN(\pipeline/stageF/PC_plus4/add_26/carry[25] ) );
  AND2_X1 \pipeline/stageF/PC_plus4/add_26/U44  ( .A1(
        \pipeline/stageF/PC_plus4/add_26/carry[23] ), .A2(addr_to_iram[23]), 
        .ZN(\pipeline/stageF/PC_plus4/add_26/carry[24] ) );
  AND2_X1 \pipeline/stageF/PC_plus4/add_26/U42  ( .A1(
        \pipeline/stageF/PC_plus4/add_26/carry[22] ), .A2(addr_to_iram[22]), 
        .ZN(\pipeline/stageF/PC_plus4/add_26/carry[23] ) );
  AND2_X1 \pipeline/stageF/PC_plus4/add_26/U40  ( .A1(
        \pipeline/stageF/PC_plus4/add_26/carry[21] ), .A2(addr_to_iram[21]), 
        .ZN(\pipeline/stageF/PC_plus4/add_26/carry[22] ) );
  AND2_X1 \pipeline/stageF/PC_plus4/add_26/U38  ( .A1(
        \pipeline/stageF/PC_plus4/add_26/carry[20] ), .A2(addr_to_iram[20]), 
        .ZN(\pipeline/stageF/PC_plus4/add_26/carry[21] ) );
  AND2_X1 \pipeline/stageF/PC_plus4/add_26/U36  ( .A1(
        \pipeline/stageF/PC_plus4/add_26/carry[19] ), .A2(addr_to_iram[19]), 
        .ZN(\pipeline/stageF/PC_plus4/add_26/carry[20] ) );
  AND2_X1 \pipeline/stageF/PC_plus4/add_26/U34  ( .A1(
        \pipeline/stageF/PC_plus4/add_26/carry[18] ), .A2(addr_to_iram[18]), 
        .ZN(\pipeline/stageF/PC_plus4/add_26/carry[19] ) );
  AND2_X1 \pipeline/stageF/PC_plus4/add_26/U32  ( .A1(
        \pipeline/stageF/PC_plus4/add_26/carry[17] ), .A2(addr_to_iram[17]), 
        .ZN(\pipeline/stageF/PC_plus4/add_26/carry[18] ) );
  AND2_X1 \pipeline/stageF/PC_plus4/add_26/U30  ( .A1(
        \pipeline/stageF/PC_plus4/add_26/carry[16] ), .A2(addr_to_iram[16]), 
        .ZN(\pipeline/stageF/PC_plus4/add_26/carry[17] ) );
  AND2_X1 \pipeline/stageF/PC_plus4/add_26/U28  ( .A1(
        \pipeline/stageF/PC_plus4/add_26/carry[15] ), .A2(addr_to_iram[15]), 
        .ZN(\pipeline/stageF/PC_plus4/add_26/carry[16] ) );
  AND2_X1 \pipeline/stageF/PC_plus4/add_26/U26  ( .A1(
        \pipeline/stageF/PC_plus4/add_26/carry[14] ), .A2(addr_to_iram[14]), 
        .ZN(\pipeline/stageF/PC_plus4/add_26/carry[15] ) );
  AND2_X1 \pipeline/stageF/PC_plus4/add_26/U24  ( .A1(
        \pipeline/stageF/PC_plus4/add_26/carry[13] ), .A2(addr_to_iram[13]), 
        .ZN(\pipeline/stageF/PC_plus4/add_26/carry[14] ) );
  AND2_X1 \pipeline/stageF/PC_plus4/add_26/U22  ( .A1(
        \pipeline/stageF/PC_plus4/add_26/carry[12] ), .A2(addr_to_iram[12]), 
        .ZN(\pipeline/stageF/PC_plus4/add_26/carry[13] ) );
  AND2_X1 \pipeline/stageF/PC_plus4/add_26/U20  ( .A1(
        \pipeline/stageF/PC_plus4/add_26/carry[11] ), .A2(addr_to_iram[11]), 
        .ZN(\pipeline/stageF/PC_plus4/add_26/carry[12] ) );
  AND2_X1 \pipeline/stageF/PC_plus4/add_26/U18  ( .A1(
        \pipeline/stageF/PC_plus4/add_26/carry[10] ), .A2(addr_to_iram[10]), 
        .ZN(\pipeline/stageF/PC_plus4/add_26/carry[11] ) );
  AND2_X1 \pipeline/stageF/PC_plus4/add_26/U16  ( .A1(
        \pipeline/stageF/PC_plus4/add_26/carry[9] ), .A2(addr_to_iram[9]), 
        .ZN(\pipeline/stageF/PC_plus4/add_26/carry[10] ) );
  AND2_X1 \pipeline/stageF/PC_plus4/add_26/U14  ( .A1(
        \pipeline/stageF/PC_plus4/add_26/carry[8] ), .A2(addr_to_iram[8]), 
        .ZN(\pipeline/stageF/PC_plus4/add_26/carry[9] ) );
  AND2_X1 \pipeline/stageF/PC_plus4/add_26/U12  ( .A1(
        \pipeline/stageF/PC_plus4/add_26/carry[7] ), .A2(addr_to_iram[7]), 
        .ZN(\pipeline/stageF/PC_plus4/add_26/carry[8] ) );
  AND2_X1 \pipeline/stageF/PC_plus4/add_26/U10  ( .A1(
        \pipeline/stageF/PC_plus4/add_26/carry[6] ), .A2(addr_to_iram[6]), 
        .ZN(\pipeline/stageF/PC_plus4/add_26/carry[7] ) );
  AND2_X1 \pipeline/stageF/PC_plus4/add_26/U8  ( .A1(
        \pipeline/stageF/PC_plus4/add_26/carry[5] ), .A2(addr_to_iram[5]), 
        .ZN(\pipeline/stageF/PC_plus4/add_26/carry[6] ) );
  AND2_X1 \pipeline/stageF/PC_plus4/add_26/U6  ( .A1(
        \pipeline/stageF/PC_plus4/add_26/carry[4] ), .A2(addr_to_iram[4]), 
        .ZN(\pipeline/stageF/PC_plus4/add_26/carry[5] ) );
  AND2_X1 \pipeline/stageF/PC_plus4/add_26/U4  ( .A1(addr_to_iram[2]), .A2(
        addr_to_iram[3]), .ZN(\pipeline/stageF/PC_plus4/add_26/carry[4] ) );
  XNOR2_X1 \pipeline/stageF/PC_plus4/add_26/U1  ( .A(addr_to_iram[30]), .B(
        \pipeline/stageF/PC_plus4/add_26/n1 ), .ZN(
        \pipeline/stageF/PC_plus4/N37 ) );
  NAND2_X1 \pipeline/stageF/PC_plus4/add_26/U2  ( .A1(
        \pipeline/stageF/PC_plus4/add_26/carry[29] ), .A2(addr_to_iram[29]), 
        .ZN(\pipeline/stageF/PC_plus4/add_26/n1 ) );
  XOR2_X1 \pipeline/stageF/PC_plus4/add_26/U55  ( .A(addr_to_iram[3]), .B(
        addr_to_iram[2]), .Z(\pipeline/stageF/PC_plus4/N10 ) );
  XOR2_X1 \pipeline/stageF/PC_plus4/add_26/U53  ( .A(addr_to_iram[4]), .B(
        \pipeline/stageF/PC_plus4/add_26/carry[4] ), .Z(
        \pipeline/stageF/PC_plus4/N11 ) );
  XOR2_X1 \pipeline/stageF/PC_plus4/add_26/U51  ( .A(addr_to_iram[5]), .B(
        \pipeline/stageF/PC_plus4/add_26/carry[5] ), .Z(
        \pipeline/stageF/PC_plus4/N12 ) );
  XOR2_X1 \pipeline/stageF/PC_plus4/add_26/U49  ( .A(addr_to_iram[6]), .B(
        \pipeline/stageF/PC_plus4/add_26/carry[6] ), .Z(
        \pipeline/stageF/PC_plus4/N13 ) );
  XOR2_X1 \pipeline/stageF/PC_plus4/add_26/U47  ( .A(addr_to_iram[7]), .B(
        \pipeline/stageF/PC_plus4/add_26/carry[7] ), .Z(
        \pipeline/stageF/PC_plus4/N14 ) );
  XOR2_X1 \pipeline/stageF/PC_plus4/add_26/U45  ( .A(addr_to_iram[8]), .B(
        \pipeline/stageF/PC_plus4/add_26/carry[8] ), .Z(
        \pipeline/stageF/PC_plus4/N15 ) );
  XOR2_X1 \pipeline/stageF/PC_plus4/add_26/U43  ( .A(addr_to_iram[9]), .B(
        \pipeline/stageF/PC_plus4/add_26/carry[9] ), .Z(
        \pipeline/stageF/PC_plus4/N16 ) );
  XOR2_X1 \pipeline/stageF/PC_plus4/add_26/U41  ( .A(addr_to_iram[10]), .B(
        \pipeline/stageF/PC_plus4/add_26/carry[10] ), .Z(
        \pipeline/stageF/PC_plus4/N17 ) );
  XOR2_X1 \pipeline/stageF/PC_plus4/add_26/U39  ( .A(addr_to_iram[11]), .B(
        \pipeline/stageF/PC_plus4/add_26/carry[11] ), .Z(
        \pipeline/stageF/PC_plus4/N18 ) );
  XOR2_X1 \pipeline/stageF/PC_plus4/add_26/U37  ( .A(addr_to_iram[12]), .B(
        \pipeline/stageF/PC_plus4/add_26/carry[12] ), .Z(
        \pipeline/stageF/PC_plus4/N19 ) );
  XOR2_X1 \pipeline/stageF/PC_plus4/add_26/U35  ( .A(addr_to_iram[13]), .B(
        \pipeline/stageF/PC_plus4/add_26/carry[13] ), .Z(
        \pipeline/stageF/PC_plus4/N20 ) );
  XOR2_X1 \pipeline/stageF/PC_plus4/add_26/U33  ( .A(addr_to_iram[14]), .B(
        \pipeline/stageF/PC_plus4/add_26/carry[14] ), .Z(
        \pipeline/stageF/PC_plus4/N21 ) );
  XOR2_X1 \pipeline/stageF/PC_plus4/add_26/U31  ( .A(addr_to_iram[15]), .B(
        \pipeline/stageF/PC_plus4/add_26/carry[15] ), .Z(
        \pipeline/stageF/PC_plus4/N22 ) );
  XOR2_X1 \pipeline/stageF/PC_plus4/add_26/U29  ( .A(addr_to_iram[16]), .B(
        \pipeline/stageF/PC_plus4/add_26/carry[16] ), .Z(
        \pipeline/stageF/PC_plus4/N23 ) );
  XOR2_X1 \pipeline/stageF/PC_plus4/add_26/U27  ( .A(addr_to_iram[17]), .B(
        \pipeline/stageF/PC_plus4/add_26/carry[17] ), .Z(
        \pipeline/stageF/PC_plus4/N24 ) );
  XOR2_X1 \pipeline/stageF/PC_plus4/add_26/U25  ( .A(addr_to_iram[18]), .B(
        \pipeline/stageF/PC_plus4/add_26/carry[18] ), .Z(
        \pipeline/stageF/PC_plus4/N25 ) );
  XOR2_X1 \pipeline/stageF/PC_plus4/add_26/U23  ( .A(addr_to_iram[19]), .B(
        \pipeline/stageF/PC_plus4/add_26/carry[19] ), .Z(
        \pipeline/stageF/PC_plus4/N26 ) );
  XOR2_X1 \pipeline/stageF/PC_plus4/add_26/U21  ( .A(addr_to_iram[20]), .B(
        \pipeline/stageF/PC_plus4/add_26/carry[20] ), .Z(
        \pipeline/stageF/PC_plus4/N27 ) );
  XOR2_X1 \pipeline/stageF/PC_plus4/add_26/U19  ( .A(addr_to_iram[21]), .B(
        \pipeline/stageF/PC_plus4/add_26/carry[21] ), .Z(
        \pipeline/stageF/PC_plus4/N28 ) );
  XOR2_X1 \pipeline/stageF/PC_plus4/add_26/U17  ( .A(addr_to_iram[22]), .B(
        \pipeline/stageF/PC_plus4/add_26/carry[22] ), .Z(
        \pipeline/stageF/PC_plus4/N29 ) );
  XOR2_X1 \pipeline/stageF/PC_plus4/add_26/U15  ( .A(addr_to_iram[23]), .B(
        \pipeline/stageF/PC_plus4/add_26/carry[23] ), .Z(
        \pipeline/stageF/PC_plus4/N30 ) );
  XOR2_X1 \pipeline/stageF/PC_plus4/add_26/U13  ( .A(addr_to_iram[24]), .B(
        \pipeline/stageF/PC_plus4/add_26/carry[24] ), .Z(
        \pipeline/stageF/PC_plus4/N31 ) );
  XOR2_X1 \pipeline/stageF/PC_plus4/add_26/U11  ( .A(addr_to_iram[25]), .B(
        \pipeline/stageF/PC_plus4/add_26/carry[25] ), .Z(
        \pipeline/stageF/PC_plus4/N32 ) );
  XOR2_X1 \pipeline/stageF/PC_plus4/add_26/U9  ( .A(addr_to_iram[26]), .B(
        \pipeline/stageF/PC_plus4/add_26/carry[26] ), .Z(
        \pipeline/stageF/PC_plus4/N33 ) );
  XOR2_X1 \pipeline/stageF/PC_plus4/add_26/U7  ( .A(addr_to_iram[27]), .B(
        \pipeline/stageF/PC_plus4/add_26/carry[27] ), .Z(
        \pipeline/stageF/PC_plus4/N34 ) );
  XOR2_X1 \pipeline/stageF/PC_plus4/add_26/U5  ( .A(addr_to_iram[28]), .B(
        \pipeline/stageF/PC_plus4/add_26/carry[28] ), .Z(
        \pipeline/stageF/PC_plus4/N35 ) );
  XOR2_X1 \pipeline/stageF/PC_plus4/add_26/U3  ( .A(addr_to_iram[29]), .B(
        \pipeline/stageF/PC_plus4/add_26/carry[29] ), .Z(
        \pipeline/stageF/PC_plus4/N36 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U97  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n109 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n108 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U92  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n45 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n23 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U85  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n115 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n30 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U162  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n152 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n151 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U91  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n64 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n29 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U29  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n83 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n82 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U86  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n99 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n9 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U93  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n4 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n35 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U112  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n60 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n114 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U45  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n24 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n112 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U44  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n25 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n111 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U165  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n133 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n132 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U89  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n107 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n106 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U11  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n40 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n8 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U26  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n88 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n87 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U107  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n90 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n89 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U104  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n102 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n101 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U111  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n103 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n75 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U94  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n14 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n39 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U12  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n5 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n43 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U87  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n134 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n17 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U168  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n162 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n161 ) );
  AND2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U95  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[3] ), .A2(n17302), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n158 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U100  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n164 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n163 ) );
  AND2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U110  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[3] ), .A2(n17081), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n84 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U7  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n58 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n52 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U5  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n56 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n51 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U10  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n53 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n48 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U6  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n2 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n46 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U40  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n115 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n5 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n59 ), .C2(n17297), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n116 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N119 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U41  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n8 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n31 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n10 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n81 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n12 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n80 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n116 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U56  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n20 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n5 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n21 ), .C2(n17297), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n22 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N112 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U57  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n8 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n23 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n10 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n24 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n12 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n25 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n22 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U48  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n4 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n5 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n6 ), .C2(n17297), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n7 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N114 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U49  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n8 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n9 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n10 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n11 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n12 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n13 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n7 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U50  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n64 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n5 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n71 ), .C2(n17737), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n148 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N115 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U51  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n8 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n30 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n10 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n31 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n12 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n81 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n148 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U60  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n14 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n5 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n15 ), .C2(n17297), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n16 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N113 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U61  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n8 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n17 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n10 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n18 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n12 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n19 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n16 ) );
  OAI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U70  ( .B1(n17112), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n110 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n60 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N121 ) );
  OAI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U71  ( .B1(n17112), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n91 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n60 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N122 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U64  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n32 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n40 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n91 ), .C2(n17737), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n92 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N106 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U65  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n12 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n9 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n43 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n93 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n10 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n35 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n92 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U172  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n46 ), .B2(n17077), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n48 ), .C2(n17102), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n98 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n93 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U173  ( .A1(n12649), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n51 ), .B1(
        \pipeline/stageE/input1_to_ALU [1]), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n52 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n98 ) );
  AOI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U96  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n13 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n73 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n11 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n1 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n108 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n91 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U98  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n105 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n72 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n84 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n74 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n109 ) );
  OAI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U76  ( .B1(n17112), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n27 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n60 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N127 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U174  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n20 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n40 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n41 ), .C2(n17297), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n42 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N108 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U175  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n12 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n24 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n43 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n44 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n10 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n23 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n42 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U176  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n46 ), .B2(n17087), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n48 ), .C2(n17088), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n50 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n44 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U177  ( .A1(
        \pipeline/stageE/input1_to_ALU [4]), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n51 ), .B1(
        \pipeline/stageE/input1_to_ALU [3]), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n52 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n50 ) );
  OAI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U149  ( .A1(n17095), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n56 ), .B1(n17089), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n58 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n54 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U62  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n26 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n40 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n61 ), .C2(n17297), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n62 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N107 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U63  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n12 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n30 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n43 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n63 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n10 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n29 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n62 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U170  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n46 ), .B2(n17102), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n48 ), .C2(n17087), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n66 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n63 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U171  ( .A1(
        \pipeline/stageE/input1_to_ALU [3]), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n51 ), .B1(n12649), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n52 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n66 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U58  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n26 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n5 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n27 ), .C2(n17737), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n28 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N111 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U59  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n8 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n29 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n10 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n30 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n12 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n31 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n28 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U163  ( .A1(
        \pipeline/stageE/input1_to_ALU [15]), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n51 ), .B1(
        \pipeline/stageE/input1_to_ALU [14]), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n52 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n152 ) );
  OAI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U155  ( .A1(n17082), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n56 ), .B1(n17085), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n58 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n154 ) );
  AOI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U28  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n80 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n73 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n81 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n1 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n82 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n27 ) );
  AOI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U30  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n84 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n85 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n86 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n83 ) );
  OAI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U146  ( .A1(n17089), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n56 ), .B1(n17088), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n58 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n67 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U52  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n32 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n5 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n33 ), .C2(n17737), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n34 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N110 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U53  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n8 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n35 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n10 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n9 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n12 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n11 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n34 ) );
  OAI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U160  ( .A1(n17085), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n56 ), .B1(n17090), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n58 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n94 ) );
  OAI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U151  ( .A1(n17088), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n56 ), .B1(n17087), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n58 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n100 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U54  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n36 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n5 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n37 ), .C2(n17297), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n38 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N109 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U55  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n8 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n39 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n10 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n17 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n12 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n18 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n38 ) );
  OAI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U84  ( .B1(n17112), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n15 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n60 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N129 ) );
  AOI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U34  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n76 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n73 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n77 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n1 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n75 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n15 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U43  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n111 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n40 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n112 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n5 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n113 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N120 ) );
  AOI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U46  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n12 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n78 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n10 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n79 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n114 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n113 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U38  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n99 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n5 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n68 ), .C2(n17737), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n118 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N118 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U39  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n8 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n11 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n10 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n13 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n12 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n74 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n118 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U137  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n46 ), .B2(n17097), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n48 ), .C2(n17118), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n127 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n11 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U138  ( .A1(
        \pipeline/stageE/input1_to_ALU [18]), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n51 ), .B1(
        \pipeline/stageE/input1_to_ALU [17]), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n52 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n127 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U166  ( .A1(
        \pipeline/stageE/input1_to_ALU [14]), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n51 ), .B1(
        \pipeline/stageE/input1_to_ALU [13]), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n52 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n133 ) );
  OAI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U72  ( .B1(n17112), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n61 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n60 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N123 ) );
  AOI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U88  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n85 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n105 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n80 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n84 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n106 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n61 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U90  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n73 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n81 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n1 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n31 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n107 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U114  ( .B1(n17097), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n56 ), .C1(n17096), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n58 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n150 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n31 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U115  ( .A1(
        \pipeline/stageE/input1_to_ALU [20]), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n2 ), .B1(
        \pipeline/stageE/input1_to_ALU [21]), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n53 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n150 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U116  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n46 ), .B2(n17117), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n48 ), .C2(n17115), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n149 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n81 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U117  ( .A1(
        \pipeline/stageE/input1_to_ALU [23]), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n51 ), .B1(
        \pipeline/stageE/input1_to_ALU [22]), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n52 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n149 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U66  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n134 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n5 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n69 ), .C2(n17297), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n135 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N117 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U67  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n8 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n18 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n10 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n19 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n12 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n77 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n135 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U68  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n45 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n5 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n70 ), .C2(n17297), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n136 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N116 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U69  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n8 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n24 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n10 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n25 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n12 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n79 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n136 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U134  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n46 ), .B2(n17079), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n48 ), .C2(n17096), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n143 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n24 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U136  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/A[16] ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n51 ), .B1(
        \pipeline/stageE/input1_to_ALU [15]), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n52 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n143 ) );
  OAI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U157  ( .A1(n17080), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n56 ), .B1(n17082), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n58 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n145 ) );
  OAI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U75  ( .B1(n17112), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n33 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n60 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N126 ) );
  AOI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U25  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n74 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n73 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n13 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n1 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n87 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n33 ) );
  AOI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U27  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n84 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n72 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n86 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n88 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U131  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n46 ), .B2(n17092), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n48 ), .C2(n17117), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n124 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n13 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U133  ( .A1(
        \pipeline/stageE/input1_to_ALU [22]), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n51 ), .B1(
        \pipeline/stageE/input1_to_ALU [21]), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n52 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n124 ) );
  OAI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U74  ( .B1(n17112), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n37 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n60 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N125 ) );
  AOI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U106  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n77 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n73 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n19 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n1 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n89 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n37 ) );
  AOI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U108  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n84 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n76 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n86 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n90 ) );
  OAI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U73  ( .B1(n17112), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n41 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n60 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N124 ) );
  AOI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U103  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n79 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n73 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n25 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n1 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n101 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n41 ) );
  AOI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U105  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n84 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n78 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n86 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n102 ) );
  NOR2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U42  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n103 ), .A2(n17081), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n86 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U123  ( .B1(n17118), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n56 ), .C1(n17097), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n58 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n140 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n25 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U124  ( .A1(
        \pipeline/stageE/input1_to_ALU [21]), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n2 ), .B1(
        \pipeline/stageE/input1_to_ALU [22]), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n53 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n140 ) );
  OAI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U78  ( .B1(n17112), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n6 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n60 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N130 ) );
  AOI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U32  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n72 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n73 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n74 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n1 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n75 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n6 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U127  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n46 ), .B2(n17078), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n48 ), .C2(n17093), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n121 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n74 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U128  ( .A1(
        \pipeline/stageE/input1_to_ALU [26]), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n51 ), .B1(
        \pipeline/stageE/input1_to_ALU [25]), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n52 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n121 ) );
  OAI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U77  ( .B1(n17112), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n21 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n60 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N128 ) );
  AOI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U31  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n78 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n73 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n79 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n1 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n75 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n21 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U125  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n46 ), .B2(n17115), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n48 ), .C2(n17086), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n139 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n79 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U126  ( .A1(
        \pipeline/stageE/input1_to_ALU [24]), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n51 ), .B1(
        \pipeline/stageE/input1_to_ALU [23]), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n52 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n139 ) );
  OAI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U79  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n71 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n60 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N131 ) );
  AOI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U33  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n85 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n73 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n80 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n1 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n75 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n71 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U143  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n46 ), .B2(n17093), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n48 ), .C2(n17094), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n153 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n80 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U144  ( .A1(
        \pipeline/stageE/input1_to_ALU [27]), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n51 ), .B1(
        \pipeline/stageE/input1_to_ALU [26]), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n52 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n153 ) );
  OAI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U80  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n70 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n60 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N132 ) );
  AOI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U35  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n78 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n1 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n117 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n70 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U141  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n46 ), .B2(n17094), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n48 ), .C2(n17083), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n144 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n78 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U142  ( .A1(
        \pipeline/stageE/input1_to_ALU [28]), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n51 ), .B1(
        \pipeline/stageE/input1_to_ALU [27]), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n52 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n144 ) );
  OAI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U83  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n69 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n60 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N133 ) );
  AOI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U37  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n76 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n1 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n117 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n69 ) );
  OAI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U81  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n68 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n60 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N134 ) );
  AOI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U17  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n72 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n1 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n117 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n68 ) );
  OAI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U24  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n58 ), .A2(n17094), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n56 ), .B2(n17083), .C1(n17303), 
        .C2(n17104), .ZN(\pipeline/stageE/EXE_ALU/alu_shift/C48/n72 ) );
  OAI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U82  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n59 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n60 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N135 ) );
  NAND2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U3  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/N136 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n60 ) );
  AOI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U36  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n85 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n1 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n117 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n59 ) );
  OAI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U109  ( .B1(n17081), .B2(
        n17104), .A(\pipeline/stageE/EXE_ALU/alu_shift/C48/n103 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n117 ) );
  NAND2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U185  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/N136 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[3] ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n103 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U178  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n36 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n40 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n110 ), .C2(n17737), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n155 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N105 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U179  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n12 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n17 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n43 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n156 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n10 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n39 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n155 ) );
  OAI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U183  ( .A1(n17090), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n56 ), .B1(n17095), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n58 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n157 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U180  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n46 ), .B2(n17091), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n48 ), .C2(n17077), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n160 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n156 ) );
  NAND2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U14  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n1 ), .A2(n17302), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n5 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U169  ( .A1(
        \pipeline/stageE/input1_to_ALU [13]), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n51 ), .B1(
        \pipeline/stageE/input1_to_ALU [12]), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n52 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n162 ) );
  AOI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U99  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n19 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n73 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n18 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n1 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n163 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n110 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U101  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n105 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n76 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n84 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n77 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n164 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U129  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n46 ), .B2(n17086), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n48 ), .C2(n17078), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n165 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n77 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U130  ( .A1(
        \pipeline/stageE/input1_to_ALU [25]), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n51 ), .B1(
        \pipeline/stageE/input1_to_ALU [24]), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n52 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n165 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U118  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n46 ), .B2(n17083), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n48 ), .C2(n17104), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n166 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n76 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U119  ( .A1(
        \pipeline/stageE/input1_to_ALU [29]), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n51 ), .B1(
        \pipeline/stageE/input1_to_ALU [28]), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n52 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n166 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U139  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n46 ), .B2(n17096), .C1(n17097), 
        .C2(\pipeline/stageE/EXE_ALU/alu_shift/C48/n48 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n167 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n18 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U140  ( .A1(
        \pipeline/stageE/input1_to_ALU [17]), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n51 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/A[16] ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n52 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n167 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U120  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n56 ), .B2(n17084), .C1(n17118), 
        .C2(\pipeline/stageE/EXE_ALU/alu_shift/C48/n58 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n169 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n19 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U122  ( .A1(
        \pipeline/stageE/input1_to_ALU [22]), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n2 ), .B1(
        \pipeline/stageE/input1_to_ALU [23]), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n53 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n169 ) );
  NAND2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U18  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n73 ), .A2(n17302), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n40 ) );
  NOR2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U2  ( .A1(n17081), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[3] ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n73 ) );
  OAI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U153  ( .A1(n17087), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n56 ), .B1(n17102), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n58 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n170 ) );
  NAND2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U16  ( .A1(n17742), .A2(
        n17303), .ZN(\pipeline/stageE/EXE_ALU/alu_shift/C48/n58 ) );
  NAND2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U9  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .A2(n17303), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n56 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C48/U148  ( .A(
        \pipeline/stageE/input1_to_ALU [30]), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/N136 ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n58 ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n85 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U114  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n4 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n130 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U76  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n48 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n128 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U77  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n81 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n127 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U47  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n40 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n121 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U62  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n33 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n95 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U50  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n31 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n117 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U59  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n42 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n102 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U56  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n50 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n107 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U53  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n16 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n113 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U105  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n73 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n72 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U113  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n104 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n84 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U65  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n20 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n88 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U97  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n169 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n168 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U5  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n12 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n56 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U108  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n162 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n161 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U36  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n154 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n153 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U187  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n85 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n45 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U40  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n144 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n143 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U184  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n77 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n37 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U33  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n140 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n139 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U176  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n170 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n98 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U178  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n64 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n28 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U6  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n53 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n17 ) );
  AND2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U99  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[3] ), .A2(n17302), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n131 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U101  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n135 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n134 ) );
  AND2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U112  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[3] ), .A2(n17081), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n74 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U181  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n58 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n11 ) );
  OAI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U94  ( .B1(n17112), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n29 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n4 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N216 ) );
  OAI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U87  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n6 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n4 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N209 ) );
  OAI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U82  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n3 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n4 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N211 ) );
  OAI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U84  ( .B1(n17112), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n61 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n4 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N212 ) );
  OAI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U95  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n5 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n4 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N210 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U75  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n127 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n12 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n128 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n53 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n129 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N218 ) );
  AOI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U78  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n15 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n82 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n19 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n83 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n130 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n129 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U46  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n121 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n53 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n112 ), .C2(n17302), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n122 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N219 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U48  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n56 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n68 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n19 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n71 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n15 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n69 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n122 ) );
  OAI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U91  ( .B1(n17112), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n112 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n4 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N203 ) );
  AOI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U42  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n75 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n1 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n109 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n112 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U61  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n95 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n53 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n7 ), .C2(n17302), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n96 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N224 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U63  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n56 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n31 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n19 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n63 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n15 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n97 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n96 ) );
  OAI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U90  ( .B1(n17112), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n10 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n4 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N205 ) );
  OAI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U89  ( .B1(n17112), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n36 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n4 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N204 ) );
  OAI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U88  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n7 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n4 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N208 ) );
  AOI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U30  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n98 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n70 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n99 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n1 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n84 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n7 ) );
  OAI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U85  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n8 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n4 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N207 ) );
  OAI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U86  ( .B1(n17112), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n9 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n4 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N206 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U73  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n45 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n53 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n5 ), .C2(n17302), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n80 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N226 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U74  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n56 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n50 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n19 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n48 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n15 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n81 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n80 ) );
  AOI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U38  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n82 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n70 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n83 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n1 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n84 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n5 ) );
  OAI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U93  ( .B1(n17112), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n13 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n4 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N217 ) );
  OAI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U92  ( .B1(n17112), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n38 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n4 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N215 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U49  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n117 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n53 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n36 ), .C2(n17302), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n118 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N220 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U51  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n56 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n63 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n19 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n97 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n15 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n99 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n118 ) );
  AOI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U43  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n98 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n1 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n109 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n36 ) );
  OAI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U81  ( .B1(n17112), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n46 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n4 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N214 ) );
  OAI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U83  ( .B1(n17112), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n54 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n4 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N213 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U58  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n102 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n53 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n8 ), .C2(n17302), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n103 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N223 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U60  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n56 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n40 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n19 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n68 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n15 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n71 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n103 ) );
  AOI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U29  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n75 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n70 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n69 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n1 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n84 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n8 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U55  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n107 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n53 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n9 ), .C2(n17302), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n108 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N222 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U57  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n56 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n48 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n19 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n81 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n15 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n83 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n108 ) );
  AOI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U45  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n82 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n1 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n109 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n9 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U52  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n113 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n53 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n10 ), .C2(n17302), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n114 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N221 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U54  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n56 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n57 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n19 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n90 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n15 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n92 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n114 ) );
  AOI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U44  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n91 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n1 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n109 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n10 ) );
  OAI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U110  ( .B1(n17119), .B2(
        n17081), .A(\pipeline/stageE/EXE_ALU/alu_shift/C86/n104 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n109 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U67  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n37 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n53 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n3 ), .C2(n17302), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n67 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N227 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U68  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n56 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n42 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n19 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n40 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n15 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n68 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n67 ) );
  AOI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U104  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n69 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n70 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n71 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n1 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n72 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n3 ) );
  AOI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U106  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n74 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n75 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n76 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n73 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U64  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n88 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n53 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n6 ), .C2(n17302), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n89 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N225 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U66  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n56 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n16 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n19 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n57 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n15 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n90 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n89 ) );
  AOI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U31  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n91 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n70 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n92 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n1 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n84 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n6 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U69  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n28 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n53 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n61 ), .C2(n17302), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n62 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N228 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U70  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n56 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n33 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n19 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n31 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n15 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n63 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n62 ) );
  AOI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U96  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n99 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n70 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n97 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n1 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n168 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n61 ) );
  AOI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U98  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n74 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n98 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n76 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n169 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U71  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n11 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n53 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n54 ), .C2(n17302), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n55 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N229 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U72  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n56 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n20 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n19 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n16 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n15 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n57 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n55 ) );
  AOI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U107  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n92 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n70 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n90 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n1 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n161 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n54 ) );
  AOI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U109  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n74 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n91 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n76 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n162 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U169  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n45 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n12 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n46 ), .C2(n17302), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n47 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N230 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U170  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n15 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n48 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n17 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n49 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n19 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n50 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n47 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U154  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n21 ), .B2(n17096), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n23 ), .C2(n17079), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n111 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n50 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U155  ( .A1(
        \pipeline/stageE/input1_to_ALU [19]), .A2(n17110), .B1(
        \pipeline/stageE/input1_to_ALU [20]), .B2(n17111), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n111 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U171  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n21 ), .B2(n17086), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n23 ), .C2(n17115), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n52 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n49 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U172  ( .A1(
        \pipeline/stageE/input1_to_ALU [27]), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n26 ), .B1(
        \pipeline/stageE/input1_to_ALU [28]), .B2(n17111), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n52 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U138  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n21 ), .B2(n17100), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n23 ), .C2(n15425), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n133 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n48 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U139  ( .A1(
        \pipeline/stageE/input1_to_ALU [15]), .A2(n17110), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/A[16] ), .B2(n17111), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n133 ) );
  AOI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U35  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n83 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n70 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n81 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n1 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n153 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n46 ) );
  AOI21_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U37  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n74 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n82 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n76 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n154 ) );
  NOR2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U111  ( .A1(n17081), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n104 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n76 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U144  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n21 ), .B2(n17091), .C1(n17103), 
        .C2(\pipeline/stageE/EXE_ALU/alu_shift/C86/n23 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n156 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n82 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U145  ( .A1(n17110), .A2(
        \pipeline/stageE/input1_to_ALU [3]), .B1(
        \pipeline/stageE/input1_to_ALU [4]), .B2(n17111), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n156 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U126  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n21 ), .B2(n17085), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n23 ), .C2(n17090), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n158 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n81 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U127  ( .A1(
        \pipeline/stageE/input1_to_ALU [11]), .A2(n17110), .B1(
        \pipeline/stageE/input1_to_ALU [12]), .B2(n17111), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n158 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U120  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n21 ), .B2(n17088), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n23 ), .C2(n17087), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n160 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n83 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U121  ( .A1(
        \pipeline/stageE/input1_to_ALU [7]), .A2(n17110), .B1(
        \pipeline/stageE/input1_to_ALU [8]), .B2(n17111), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n160 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U188  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n21 ), .B2(n17116), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n23 ), .C2(n17084), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n87 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n85 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U189  ( .A1(
        \pipeline/stageE/input1_to_ALU [23]), .A2(n17110), .B1(n17158), .B2(
        n17111), .ZN(\pipeline/stageE/EXE_ALU/alu_shift/C86/n87 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U156  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n37 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n12 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n38 ), .C2(n17302), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n39 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N231 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U157  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n15 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n40 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n17 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n41 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n19 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n42 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n39 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U148  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n21 ), .B2(n17097), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n23 ), .C2(n17096), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n106 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n42 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U149  ( .A1(
        \pipeline/stageE/input1_to_ALU [20]), .A2(n17110), .B1(
        \pipeline/stageE/input1_to_ALU [21]), .B2(n17111), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n106 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U158  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n21 ), .B2(n17078), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n23 ), .C2(n17086), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n44 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n41 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U159  ( .A1(
        \pipeline/stageE/input1_to_ALU [28]), .A2(n17110), .B1(
        \pipeline/stageE/input1_to_ALU [29]), .B2(n17111), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n44 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U132  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n21 ), .B2(n17101), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n23 ), .C2(n17100), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n126 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n40 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U133  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/A[16] ), .A2(n17110), .B1(
        \pipeline/stageE/input1_to_ALU [17]), .B2(n17111), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n126 ) );
  AOI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U39  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n75 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n136 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n69 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n74 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n143 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n38 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U41  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n70 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n71 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n1 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n68 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n144 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U174  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n21 ), .B2(n17082), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n23 ), .C2(n17085), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n146 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n68 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U175  ( .A1(
        \pipeline/stageE/input1_to_ALU [12]), .A2(n17110), .B1(
        \pipeline/stageE/input1_to_ALU [13]), .B2(n17111), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n146 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U116  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n21 ), .B2(n17089), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n23 ), .C2(n17088), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n149 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n71 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U117  ( .A1(
        \pipeline/stageE/input1_to_ALU [8]), .A2(n17110), .B1(
        \pipeline/stageE/input1_to_ALU [9]), .B2(n17111), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n149 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U146  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n21 ), .B2(n17077), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n23 ), .C2(n17091), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n152 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n69 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U147  ( .A1(
        \pipeline/stageE/input1_to_ALU [4]), .A2(n17110), .B1(
        \pipeline/stageE/input1_to_ALU [5]), .B2(n17111), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n152 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U185  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n21 ), .B2(n17092), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n23 ), .C2(n17116), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n79 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n77 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U186  ( .A1(n17158), .A2(
        n17110), .B1(n17159), .B2(n17111), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n79 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U160  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n28 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n12 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n29 ), .C2(n17302), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n30 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N232 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U161  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n15 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n31 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n17 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n32 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n19 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n33 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n30 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U150  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n21 ), .B2(n17118), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n23 ), .C2(n17097), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n101 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n33 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U151  ( .A1(
        \pipeline/stageE/input1_to_ALU [21]), .A2(n17110), .B1(
        \pipeline/stageE/input1_to_ALU [22]), .B2(n17111), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n101 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U162  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n21 ), .B2(n17093), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n23 ), .C2(n17078), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n35 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n32 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U163  ( .A1(
        \pipeline/stageE/input1_to_ALU [29]), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n26 ), .B1(
        \pipeline/stageE/input1_to_ALU [30]), .B2(n17111), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n35 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U134  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n21 ), .B2(n17738), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n23 ), .C2(n17101), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n120 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n31 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U135  ( .A1(
        \pipeline/stageE/input1_to_ALU [17]), .A2(n17110), .B1(
        \pipeline/stageE/input1_to_ALU [18]), .B2(n17111), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n120 ) );
  AOI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U32  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n97 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n70 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n63 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n1 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n139 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n29 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U34  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n136 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n98 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n74 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n99 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n140 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U122  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n21 ), .B2(n17102), .C1(n17077), 
        .C2(\pipeline/stageE/EXE_ALU/alu_shift/C86/n23 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n172 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n99 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U123  ( .A1(
        \pipeline/stageE/input1_to_ALU [5]), .A2(n17110), .B1(
        \pipeline/stageE/input1_to_ALU [6]), .B2(n17111), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n172 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U140  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n21 ), .B2(n17080), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n23 ), .C2(n17082), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n142 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n63 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U141  ( .A1(n17160), .A2(
        n17110), .B1(\pipeline/stageE/input1_to_ALU [14]), .B2(n17111), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n142 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U128  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n21 ), .B2(n17095), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n23 ), .C2(n17089), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n171 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n97 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U129  ( .A1(
        \pipeline/stageE/input1_to_ALU [9]), .A2(n17110), .B1(
        \pipeline/stageE/input1_to_ALU [10]), .B2(n17111), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n171 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U179  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n21 ), .B2(n17117), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n23 ), .C2(n17092), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n66 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n64 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U180  ( .A1(n17159), .A2(
        n17110), .B1(\pipeline/stageE/input1_to_ALU [26]), .B2(n17111), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n66 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U164  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n11 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n12 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n13 ), .C2(n17302), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n14 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N233 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U166  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n15 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n16 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n17 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n18 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n19 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n20 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n14 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U152  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n21 ), .B2(n17084), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n23 ), .C2(n17118), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n94 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n20 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U153  ( .A1(
        \pipeline/stageE/input1_to_ALU [22]), .A2(n17110), .B1(
        \pipeline/stageE/input1_to_ALU [23]), .B2(n17111), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n94 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U167  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n21 ), .B2(n17094), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n23 ), .C2(n17093), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n25 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n18 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U173  ( .A1(
        \pipeline/stageE/input1_to_ALU [30]), .A2(n17110), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/N136 ), .B2(n17111), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n25 ) );
  NAND2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U14  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n1 ), .A2(n17302), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n53 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U136  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n21 ), .B2(n17079), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n23 ), .C2(n17738), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n116 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n16 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U137  ( .A1(
        \pipeline/stageE/input1_to_ALU [18]), .A2(n17110), .B1(
        \pipeline/stageE/input1_to_ALU [19]), .B2(n17111), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n116 ) );
  AOI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U100  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n90 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n70 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n57 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n1 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n134 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n13 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U102  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n136 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n91 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n74 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n92 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n135 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U124  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n21 ), .B2(n17087), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n23 ), .C2(n17102), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n167 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n92 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U125  ( .A1(
        \pipeline/stageE/input1_to_ALU [6]), .A2(n17110), .B1(
        \pipeline/stageE/input1_to_ALU [7]), .B2(n17111), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n167 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U118  ( .B1(n17103), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n21 ), .C1(n17119), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n23 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n163 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n91 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U119  ( .A1(n17110), .A2(
        n12649), .B1(\pipeline/stageE/input1_to_ALU [3]), .B2(n17111), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n163 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U142  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n21 ), .B2(n15425), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n23 ), .C2(n17080), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n138 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n57 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U143  ( .A1(
        \pipeline/stageE/input1_to_ALU [14]), .A2(n17110), .B1(
        \pipeline/stageE/input1_to_ALU [15]), .B2(n17111), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n138 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U130  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n21 ), .B2(n17090), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n23 ), .C2(n17095), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n165 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n90 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U131  ( .A1(
        \pipeline/stageE/input1_to_ALU [10]), .A2(n17110), .B1(
        \pipeline/stageE/input1_to_ALU [11]), .B2(n17111), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n165 ) );
  NAND2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U15  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n70 ), .A2(n17302), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n12 ) );
  NOR2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U2  ( .A1(n17081), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[3] ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n70 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U182  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n21 ), .B2(n17115), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n23 ), .C2(n17117), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n60 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n58 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U183  ( .A1(
        \pipeline/stageE/input1_to_ALU [26]), .A2(n17110), .B1(
        \pipeline/stageE/input1_to_ALU [27]), .B2(n17111), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n60 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C86/U165  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/N202 ), .B(
        \pipeline/stageE/input1_to_ALU [1]), .S(n17111), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n75 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M0_0_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/N202 ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/N136 ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][0] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_0_1  ( .A(
        \pipeline/stageE/input1_to_ALU [1]), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/N202 ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][1] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_0_2  ( .A(n12649), .B(
        \pipeline/stageE/input1_to_ALU [1]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][2] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_0_3  ( .A(
        \pipeline/stageE/input1_to_ALU [3]), .B(n12649), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][3] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_0_5  ( .A(
        \pipeline/stageE/input1_to_ALU [5]), .B(
        \pipeline/stageE/input1_to_ALU [4]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][5] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_0_6  ( .A(
        \pipeline/stageE/input1_to_ALU [6]), .B(
        \pipeline/stageE/input1_to_ALU [5]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][6] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_0_7  ( .A(
        \pipeline/stageE/input1_to_ALU [7]), .B(
        \pipeline/stageE/input1_to_ALU [6]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][7] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_0_8  ( .A(
        \pipeline/stageE/input1_to_ALU [8]), .B(
        \pipeline/stageE/input1_to_ALU [7]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][8] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_0_9  ( .A(
        \pipeline/stageE/input1_to_ALU [9]), .B(
        \pipeline/stageE/input1_to_ALU [8]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][9] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_0_10  ( .A(
        \pipeline/stageE/input1_to_ALU [10]), .B(
        \pipeline/stageE/input1_to_ALU [9]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][10] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_0_11  ( .A(
        \pipeline/stageE/input1_to_ALU [11]), .B(
        \pipeline/stageE/input1_to_ALU [10]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][11] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_0_12  ( .A(
        \pipeline/stageE/input1_to_ALU [12]), .B(
        \pipeline/stageE/input1_to_ALU [11]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][12] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_0_13  ( .A(
        \pipeline/stageE/input1_to_ALU [13]), .B(
        \pipeline/stageE/input1_to_ALU [12]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][13] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_0_14  ( .A(
        \pipeline/stageE/input1_to_ALU [14]), .B(
        \pipeline/stageE/input1_to_ALU [13]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][14] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_0_15  ( .A(
        \pipeline/stageE/input1_to_ALU [15]), .B(
        \pipeline/stageE/input1_to_ALU [14]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][15] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_0_16  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/A[16] ), .B(
        \pipeline/stageE/input1_to_ALU [15]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][16] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_0_17  ( .A(
        \pipeline/stageE/input1_to_ALU [17]), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/A[16] ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][17] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_0_18  ( .A(
        \pipeline/stageE/input1_to_ALU [18]), .B(
        \pipeline/stageE/input1_to_ALU [17]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][18] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_0_19  ( .A(
        \pipeline/stageE/input1_to_ALU [19]), .B(
        \pipeline/stageE/input1_to_ALU [18]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][19] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_0_20  ( .A(
        \pipeline/stageE/input1_to_ALU [20]), .B(
        \pipeline/stageE/input1_to_ALU [19]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][20] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_0_21  ( .A(
        \pipeline/stageE/input1_to_ALU [21]), .B(
        \pipeline/stageE/input1_to_ALU [20]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][21] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_0_22  ( .A(
        \pipeline/stageE/input1_to_ALU [22]), .B(
        \pipeline/stageE/input1_to_ALU [21]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][22] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_0_23  ( .A(
        \pipeline/stageE/input1_to_ALU [23]), .B(
        \pipeline/stageE/input1_to_ALU [22]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][23] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_0_24  ( .A(
        \pipeline/stageE/input1_to_ALU [24]), .B(
        \pipeline/stageE/input1_to_ALU [23]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][24] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_0_25  ( .A(
        \pipeline/stageE/input1_to_ALU [25]), .B(
        \pipeline/stageE/input1_to_ALU [24]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][25] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_0_26  ( .A(
        \pipeline/stageE/input1_to_ALU [26]), .B(
        \pipeline/stageE/input1_to_ALU [25]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][26] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_0_27  ( .A(
        \pipeline/stageE/input1_to_ALU [27]), .B(
        \pipeline/stageE/input1_to_ALU [26]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][27] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_0_28  ( .A(
        \pipeline/stageE/input1_to_ALU [28]), .B(
        \pipeline/stageE/input1_to_ALU [27]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][28] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_0_29  ( .A(
        \pipeline/stageE/input1_to_ALU [29]), .B(
        \pipeline/stageE/input1_to_ALU [28]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][29] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_0_30  ( .A(
        \pipeline/stageE/input1_to_ALU [30]), .B(
        \pipeline/stageE/input1_to_ALU [29]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][30] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_0_31  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/N136 ), .B(
        \pipeline/stageE/input1_to_ALU [30]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][31] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M0_1_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][0] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][30] ), .S(n17099), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][0] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M0_1_1  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][1] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][31] ), .S(n17099), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][1] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_1_2  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][2] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][0] ), .S(n17099), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][2] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_1_3  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][3] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][1] ), .S(n17298), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][3] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_1_4  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][4] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][2] ), .S(n17099), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][4] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_1_5  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][5] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][3] ), .S(n17298), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][5] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_1_6  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][6] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][4] ), .S(n17298), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][6] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_1_7  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][7] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][5] ), .S(n17298), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][7] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_1_8  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][8] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][6] ), .S(n17099), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][8] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_1_9  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][9] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][7] ), .S(n17298), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][9] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_1_10  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][10] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][8] ), .S(n17099), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][10] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_1_11  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][11] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][9] ), .S(n17099), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][11] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_1_12  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][12] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][10] ), .S(n17099), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][12] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_1_13  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][13] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][11] ), .S(n17298), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][13] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_1_14  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][14] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][12] ), .S(n17099), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][14] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_1_15  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][15] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][13] ), .S(n17099), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][15] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_1_16  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][16] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][14] ), .S(n17298), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][16] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_1_17  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][17] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][15] ), .S(n17099), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][17] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_1_18  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][18] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][16] ), .S(n17099), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][18] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_1_19  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][19] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][17] ), .S(n17298), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][19] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_1_20  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][20] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][18] ), .S(n17298), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][20] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_1_21  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][21] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][19] ), .S(n17099), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][21] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_1_22  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][22] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][20] ), .S(n17099), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][22] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_1_23  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][23] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][21] ), .S(n17099), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][23] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_1_24  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][24] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][22] ), .S(n17099), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][24] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_1_25  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][25] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][23] ), .S(n17298), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][25] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_1_26  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][26] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][24] ), .S(n17099), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][26] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_1_27  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][27] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][25] ), .S(n17298), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][27] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_1_28  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][28] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][26] ), .S(n17099), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][28] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_1_29  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][29] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][27] ), .S(n17099), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][29] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_1_30  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][30] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][28] ), .S(n17099), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][30] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_1_31  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][31] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[1][29] ), .S(n17099), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][31] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M0_2_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][0] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][28] ), .S(n17114), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][0] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M0_2_1  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][1] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][29] ), .S(n17114), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][1] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M0_2_2  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][2] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][30] ), .S(n17114), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][2] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M0_2_3  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][3] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][31] ), .S(n17114), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][3] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_2_4  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][4] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][0] ), .S(n17074), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][4] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_2_5  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][5] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][1] ), .S(n17114), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][5] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_2_6  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][6] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][2] ), .S(n17074), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][6] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_2_7  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][7] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][3] ), .S(n17114), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][7] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_2_8  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][8] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][4] ), .S(n17074), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][8] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_2_9  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][9] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][5] ), .S(n17074), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][9] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_2_10  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][10] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][6] ), .S(n17074), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][10] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_2_11  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][11] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][7] ), .S(n17074), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][11] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_2_12  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][12] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][8] ), .S(n17074), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][12] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_2_13  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][13] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][9] ), .S(n17074), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][13] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_2_14  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][14] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][10] ), .S(n17114), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][14] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_2_15  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][15] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][11] ), .S(n17114), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][15] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_2_16  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][16] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][12] ), .S(n17074), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][16] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_2_17  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][17] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][13] ), .S(n17114), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][17] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_2_18  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][18] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][14] ), .S(n17114), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][18] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_2_19  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][19] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][15] ), .S(n17114), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][19] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_2_20  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][20] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][16] ), .S(n17114), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][20] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_2_21  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][21] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][17] ), .S(n17114), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][21] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_2_22  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][22] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][18] ), .S(n17074), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][22] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_2_23  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][23] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][19] ), .S(n17074), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][23] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_2_24  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][24] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][20] ), .S(n17074), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][24] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_2_25  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][25] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][21] ), .S(n17074), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][25] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_2_26  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][26] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][22] ), .S(n17074), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][26] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_2_27  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][27] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][23] ), .S(n17074), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][27] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_2_28  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][28] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][24] ), .S(n17074), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][28] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_2_29  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][29] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][25] ), .S(n17074), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][29] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_2_30  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][30] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][26] ), .S(n17074), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][30] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_2_31  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][31] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[2][27] ), .S(n17074), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][31] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M0_3_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][0] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][24] ), .S(n17301), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][0] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M0_3_1  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][1] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][25] ), .S(n17301), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][1] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M0_3_2  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][2] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][26] ), .S(n17301), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][2] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M0_3_3  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][3] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][27] ), .S(n17301), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][3] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M0_3_4  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][4] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][28] ), .S(n17301), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][4] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M0_3_5  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][5] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][29] ), .S(n17301), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][5] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M0_3_6  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][6] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][30] ), .S(n17301), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][6] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M0_3_7  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][7] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][31] ), .S(n17301), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][7] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_3_8  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][8] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][0] ), .S(n17301), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][8] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_3_9  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][9] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][1] ), .S(n17301), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][9] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_3_10  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][10] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][2] ), .S(n17301), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][10] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_3_11  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][11] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][3] ), .S(n17301), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][11] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_3_12  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][12] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][4] ), .S(n17300), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][12] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_3_13  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][13] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][5] ), .S(n17300), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][13] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_3_14  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][14] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][6] ), .S(n17300), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][14] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_3_15  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][15] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][7] ), .S(n17300), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][15] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_3_16  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][16] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][8] ), .S(n17300), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][16] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_3_17  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][17] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][9] ), .S(n17300), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][17] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_3_18  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][18] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][10] ), .S(n17300), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][18] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_3_19  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][19] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][11] ), .S(n17300), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][19] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_3_20  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][20] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][12] ), .S(n17300), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][20] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_3_21  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][21] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][13] ), .S(n17300), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][21] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_3_22  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][22] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][14] ), .S(n17300), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][22] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_3_23  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][23] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][15] ), .S(n17300), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][23] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_3_24  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][24] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][16] ), .S(n17301), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][24] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_3_25  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][25] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][17] ), .S(n17300), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][25] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_3_26  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][26] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][18] ), .S(n17300), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][26] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_3_27  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][27] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][19] ), .S(n17299), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][27] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_3_28  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][28] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][20] ), .S(n17299), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][28] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_3_29  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][29] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][21] ), .S(n17299), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][29] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_3_30  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][30] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][22] ), .S(n17299), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][30] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_3_31  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][31] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[3][23] ), .S(n17300), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][31] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M0_4_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][0] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][16] ), .S(n17112), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/N39 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M0_4_1  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][1] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][17] ), .S(n17112), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/N40 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M0_4_2  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][2] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][18] ), .S(n17112), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/N41 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M0_4_3  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][3] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][19] ), .S(n17112), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/N42 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M0_4_4  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][4] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][20] ), .S(n17112), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/N43 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M0_4_5  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][5] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][21] ), .S(n17112), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/N44 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M0_4_6  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][6] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][22] ), .S(n17112), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/N45 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M0_4_7  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][7] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][23] ), .S(n17112), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/N46 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M0_4_8  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][8] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][24] ), .S(n17112), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/N47 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M0_4_9  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][9] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][25] ), .S(n17112), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/N48 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M0_4_10  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][10] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][26] ), .S(n17112), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/N49 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M0_4_11  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][11] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][27] ), .S(n17112), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/N50 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M0_4_12  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][12] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][28] ), .S(n17112), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/N51 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M0_4_13  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][13] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][29] ), .S(n17112), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/N52 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M0_4_14  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][14] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][30] ), .S(n17112), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/N53 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M0_4_15  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][15] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][31] ), .S(n17112), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/N54 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_4_16  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][16] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][0] ), .S(n17112), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N55 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_4_17  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][17] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][1] ), .S(n17112), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N56 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_4_18  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][18] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][2] ), .S(n17112), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N57 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_4_19  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][19] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][3] ), .S(n17112), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N58 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_4_20  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][20] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][4] ), .S(n17112), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N59 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_4_21  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][21] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][5] ), .S(n17112), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N60 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_4_22  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][22] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][6] ), .S(n17112), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N61 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_4_23  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][23] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][7] ), .S(n17112), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N62 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_4_24  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][24] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][8] ), .S(n17112), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N63 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_4_25  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][25] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][9] ), .S(n17112), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N64 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_4_26  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][26] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][10] ), .S(n17112), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/N65 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_4_27  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][27] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][11] ), .S(n17112), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/N66 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_4_28  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][28] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][12] ), .S(n17112), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/N67 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_4_29  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][29] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][13] ), .S(n17112), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/N68 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_4_30  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][30] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][14] ), .S(n17112), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/N69 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C10/M1_4_31  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][31] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C10/ML_int[4][15] ), .S(n17112), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/N70 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_0_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/N202 ), .B(
        \pipeline/stageE/input1_to_ALU [1]), .S(n17113), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][0] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_0_1_0  ( .A(
        \pipeline/stageE/input1_to_ALU [1]), .B(n12649), .S(n17113), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][1] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_0_2_0  ( .A(n12649), .B(
        \pipeline/stageE/input1_to_ALU [3]), .S(n17113), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][2] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_0_3_0  ( .A(
        \pipeline/stageE/input1_to_ALU [3]), .B(
        \pipeline/stageE/input1_to_ALU [4]), .S(n17113), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][3] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_0_4_0  ( .A(
        \pipeline/stageE/input1_to_ALU [4]), .B(
        \pipeline/stageE/input1_to_ALU [5]), .S(n17113), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][4] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_0_5_0  ( .A(
        \pipeline/stageE/input1_to_ALU [5]), .B(
        \pipeline/stageE/input1_to_ALU [6]), .S(n17113), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][5] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_0_6_0  ( .A(
        \pipeline/stageE/input1_to_ALU [6]), .B(
        \pipeline/stageE/input1_to_ALU [7]), .S(n17113), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][6] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_0_7_0  ( .A(
        \pipeline/stageE/input1_to_ALU [7]), .B(
        \pipeline/stageE/input1_to_ALU [8]), .S(n17113), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][7] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_0_8_0  ( .A(
        \pipeline/stageE/input1_to_ALU [8]), .B(
        \pipeline/stageE/input1_to_ALU [9]), .S(n17113), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][8] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_0_9_0  ( .A(
        \pipeline/stageE/input1_to_ALU [9]), .B(
        \pipeline/stageE/input1_to_ALU [10]), .S(n17113), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][9] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_0_10_0  ( .A(
        \pipeline/stageE/input1_to_ALU [10]), .B(
        \pipeline/stageE/input1_to_ALU [11]), .S(n17113), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][10] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_0_11_0  ( .A(
        \pipeline/stageE/input1_to_ALU [11]), .B(
        \pipeline/stageE/input1_to_ALU [12]), .S(n17113), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][11] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_0_12_0  ( .A(
        \pipeline/stageE/input1_to_ALU [12]), .B(
        \pipeline/stageE/input1_to_ALU [13]), .S(n17113), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][12] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_0_13_0  ( .A(
        \pipeline/stageE/input1_to_ALU [13]), .B(
        \pipeline/stageE/input1_to_ALU [14]), .S(n17113), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][13] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_0_14_0  ( .A(
        \pipeline/stageE/input1_to_ALU [14]), .B(
        \pipeline/stageE/input1_to_ALU [15]), .S(n17113), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][14] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_0_15_0  ( .A(
        \pipeline/stageE/input1_to_ALU [15]), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/A[16] ), .S(n17113), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][15] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_0_16_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/A[16] ), .B(
        \pipeline/stageE/input1_to_ALU [17]), .S(n17113), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][16] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_0_17_0  ( .A(
        \pipeline/stageE/input1_to_ALU [17]), .B(
        \pipeline/stageE/input1_to_ALU [18]), .S(n17113), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][17] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_0_18_0  ( .A(
        \pipeline/stageE/input1_to_ALU [18]), .B(
        \pipeline/stageE/input1_to_ALU [19]), .S(n17113), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][18] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_0_19_0  ( .A(
        \pipeline/stageE/input1_to_ALU [19]), .B(
        \pipeline/stageE/input1_to_ALU [20]), .S(n17113), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][19] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_0_20_0  ( .A(
        \pipeline/stageE/input1_to_ALU [20]), .B(
        \pipeline/stageE/input1_to_ALU [21]), .S(n17113), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][20] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_0_21_0  ( .A(
        \pipeline/stageE/input1_to_ALU [21]), .B(
        \pipeline/stageE/input1_to_ALU [22]), .S(n17113), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][21] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_0_22_0  ( .A(
        \pipeline/stageE/input1_to_ALU [22]), .B(
        \pipeline/stageE/input1_to_ALU [23]), .S(n17113), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][22] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_0_23_0  ( .A(
        \pipeline/stageE/input1_to_ALU [23]), .B(
        \pipeline/stageE/input1_to_ALU [24]), .S(n17113), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][23] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_0_24_0  ( .A(
        \pipeline/stageE/input1_to_ALU [24]), .B(
        \pipeline/stageE/input1_to_ALU [25]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][24] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_0_25_0  ( .A(
        \pipeline/stageE/input1_to_ALU [25]), .B(
        \pipeline/stageE/input1_to_ALU [26]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][25] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_0_26_0  ( .A(
        \pipeline/stageE/input1_to_ALU [26]), .B(
        \pipeline/stageE/input1_to_ALU [27]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][26] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_0_27_0  ( .A(
        \pipeline/stageE/input1_to_ALU [27]), .B(
        \pipeline/stageE/input1_to_ALU [28]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][27] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_0_28_0  ( .A(
        \pipeline/stageE/input1_to_ALU [28]), .B(
        \pipeline/stageE/input1_to_ALU [29]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][28] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_0_29_0  ( .A(
        \pipeline/stageE/input1_to_ALU [29]), .B(
        \pipeline/stageE/input1_to_ALU [30]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][29] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_0_30_0  ( .A(
        \pipeline/stageE/input1_to_ALU [30]), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/N136 ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][30] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_0_31_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/N136 ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/N202 ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][31] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_1_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][0] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][2] ), .S(n17099), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][0] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_1_1  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][1] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][3] ), .S(n17099), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][1] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_1_2_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][2] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][4] ), .S(n17099), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][2] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_1_3_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][3] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][5] ), .S(n17099), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][3] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_1_4_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][4] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][6] ), .S(n17099), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][4] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_1_5_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][5] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][7] ), .S(n17099), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][5] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_1_6_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][6] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][8] ), .S(n17099), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][6] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_1_7_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][7] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][9] ), .S(n17099), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][7] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_1_8_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][8] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][10] ), .S(n17099), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][8] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_1_9_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][9] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][11] ), .S(n17099), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][9] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_1_10_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][10] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][12] ), .S(n17099), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][10] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_1_11_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][11] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][13] ), .S(n17099), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][11] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_1_12_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][12] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][14] ), .S(n17298), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][12] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_1_13_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][13] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][15] ), .S(n17298), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][13] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_1_14_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][14] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][16] ), .S(n17298), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][14] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_1_15_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][15] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][17] ), .S(n17298), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][15] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_1_16_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][16] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][18] ), .S(n17298), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][16] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_1_17_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][17] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][19] ), .S(n17298), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][17] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_1_18_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][18] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][20] ), .S(n17298), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][18] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_1_19_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][19] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][21] ), .S(n17298), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][19] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_1_20_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][20] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][22] ), .S(n17298), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][20] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_1_21_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][21] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][23] ), .S(n17298), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][21] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_1_22_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][22] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][24] ), .S(n17298), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][22] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_1_23_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][23] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][25] ), .S(n17298), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][23] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_1_24_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][24] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][26] ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[1] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][24] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_1_25_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][25] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][27] ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[1] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][25] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_1_26_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][26] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][28] ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[1] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][26] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_1_27_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][27] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][29] ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[1] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][27] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_1_28_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][28] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][30] ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[1] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][28] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_1_29_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][29] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][31] ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[1] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][29] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_1_30_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][30] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][0] ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[1] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][30] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_1_31_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][31] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[1][1] ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[1] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][31] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_2_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][0] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][4] ), .S(n17074), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][0] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_2_1  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][1] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][5] ), .S(n17074), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][1] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_2_2  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][2] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][6] ), .S(n17074), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][2] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_2_3  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][3] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][7] ), .S(n17114), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][3] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_2_4_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][4] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][8] ), .S(n17114), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][4] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_2_5_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][5] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][9] ), .S(n17074), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][5] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_2_6_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][6] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][10] ), .S(n17074), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][6] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_2_7_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][7] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][11] ), .S(n17114), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][7] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_2_8_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][8] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][12] ), .S(n17114), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][8] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_2_9_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][9] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][13] ), .S(n17074), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][9] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_2_10_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][10] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][14] ), .S(n17074), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][10] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_2_11_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][11] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][15] ), .S(n17074), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][11] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_2_12_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][12] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][16] ), .S(n17074), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][12] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_2_13_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][13] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][17] ), .S(n17074), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][13] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_2_14_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][14] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][18] ), .S(n17074), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][14] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_2_15_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][15] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][19] ), .S(n17074), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][15] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_2_16_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][16] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][20] ), .S(n17074), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][16] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_2_17_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][17] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][21] ), .S(n17074), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][17] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_2_18_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][18] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][22] ), .S(n17074), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][18] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_2_19_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][19] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][23] ), .S(n17074), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][19] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_2_20_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][20] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][24] ), .S(n17074), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][20] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_2_21_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][21] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][25] ), .S(n17074), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][21] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_2_22_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][22] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][26] ), .S(n17074), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][22] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_2_23_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][23] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][27] ), .S(n17074), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][23] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_2_24_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][24] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][28] ), .S(n17074), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][24] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_2_25_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][25] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][29] ), .S(n17074), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][25] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_2_26_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][26] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][30] ), .S(n17074), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][26] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_2_27_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][27] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][31] ), .S(n17074), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][27] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_2_28_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][28] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][0] ), .S(n17074), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][28] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_2_29_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][29] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][1] ), .S(n17074), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][29] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_2_30_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][30] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][2] ), .S(n17074), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][30] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_2_31_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][31] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[2][3] ), .S(n17074), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][31] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_3_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][0] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][8] ), .S(n17299), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][0] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_3_1  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][1] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][9] ), .S(n17299), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][1] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_3_2  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][2] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][10] ), .S(n17299), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][2] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_3_3  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][3] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][11] ), .S(n17299), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][3] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_3_4  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][4] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][12] ), .S(n17299), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][4] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_3_5  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][5] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][13] ), .S(n17299), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][5] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_3_6  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][6] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][14] ), .S(n17299), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][6] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_3_7  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][7] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][15] ), .S(n17299), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][7] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_3_8_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][8] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][16] ), .S(n17299), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][8] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_3_9_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][9] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][17] ), .S(n17299), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][9] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_3_10_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][10] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][18] ), .S(n17299), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][10] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_3_11_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][11] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][19] ), .S(n17299), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][11] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_3_12_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][12] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][20] ), .S(n17296), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][12] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_3_13_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][13] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][21] ), .S(n17296), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][13] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_3_14_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][14] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][22] ), .S(n17296), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][14] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_3_15_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][15] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][23] ), .S(n17296), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][15] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_3_16_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][16] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][24] ), .S(n17296), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][16] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_3_17_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][17] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][25] ), .S(n17296), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][17] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_3_18_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][18] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][26] ), .S(n17296), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][18] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_3_19_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][19] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][27] ), .S(n17296), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][19] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_3_20_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][20] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][28] ), .S(n17296), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][20] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_3_21_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][21] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][29] ), .S(n17296), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][21] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_3_22_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][22] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][30] ), .S(n17296), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][22] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_3_23_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][23] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][31] ), .S(n17296), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][23] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_3_24_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][24] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][0] ), .S(n17300), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][24] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_3_25_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][25] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][1] ), .S(n17299), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][25] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_3_26_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][26] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][2] ), .S(n17301), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][26] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_3_27_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][27] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][3] ), .S(n17301), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][27] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_3_28_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][28] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][4] ), .S(n17296), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][28] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_3_29_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][29] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][5] ), .S(n17296), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][29] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_3_30_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][30] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][6] ), .S(n17301), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][30] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_3_31_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][31] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[3][7] ), .S(n17299), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][31] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_4_0  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][0] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][16] ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N7 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_4_1  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][1] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][17] ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N8 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_4_2  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][2] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][18] ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N9 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_4_3  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][3] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][19] ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N10 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_4_4  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][4] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][20] ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N11 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_4_5  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][5] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][21] ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N12 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_4_6  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][6] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][22] ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N13 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_4_7  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][7] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][23] ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N14 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_4_8  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][8] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][24] ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N15 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_4_9  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][9] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][25] ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N16 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_4_10  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][10] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][26] ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N17 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_4_11  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][11] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][27] ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N18 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_4_12  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][12] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][28] ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N19 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_4_13  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][13] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][29] ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N20 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_4_14  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][14] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][30] ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N21 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_4_15  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][15] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][31] ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N22 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_4_16  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][16] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][0] ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N23 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_4_17  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][17] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][1] ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N24 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_4_18  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][18] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][2] ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N25 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_4_19  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][19] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][3] ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N26 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_4_20  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][20] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][4] ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N27 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_4_21  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][21] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][5] ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N28 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_4_22  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][22] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][6] ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N29 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_4_23  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][23] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][7] ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N30 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_4_24  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][24] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][8] ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N31 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_4_25  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][25] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][9] ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N32 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_4_26  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][26] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][10] ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N33 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_4_27  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][27] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][11] ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N34 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_4_28  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][28] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][12] ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N35 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_4_29  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][29] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][13] ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N36 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_4_30  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][30] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][14] ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N37 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C8/M1_4_31  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][31] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C8/MR_int[4][15] ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N38 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U87  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n28 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n101 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U88  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n29 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n100 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U107  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n94 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n93 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U100  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n43 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n21 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U96  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n63 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n27 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U97  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n2 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n33 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U84  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n23 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n96 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U80  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n7 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n104 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U81  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n9 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n103 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U110  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n91 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n90 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U101  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n121 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N149 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U104  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n123 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n122 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U8  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n38 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n6 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U99  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n22 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n97 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U44  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n89 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n69 ) );
  AND2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U112  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n68 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n41 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N165 ) );
  AND2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U46  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n67 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n41 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N166 ) );
  AND2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U47  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n59 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n41 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N167 ) );
  AND2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U48  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n41 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n58 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N168 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U98  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n12 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n37 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U5  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n3 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n41 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U59  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n156 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n155 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U9  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n50 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n57 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U7  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n49 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n55 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U11  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n44 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n51 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U86  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n100 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n38 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n101 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n3 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n102 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N151 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U89  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n10 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n78 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n99 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n59 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n8 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n79 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n102 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U70  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n18 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n3 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n19 ), .C2(n17297), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n20 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N144 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U71  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n6 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n21 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n8 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n22 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n10 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n23 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n20 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U62  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n2 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n3 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n4 ), .C2(n17297), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n5 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N146 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U63  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n6 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n7 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n8 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n9 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n10 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n11 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n5 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U64  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n63 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n3 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n70 ), .C2(n17297), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n138 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N147 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U65  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n6 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n28 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n8 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n29 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n10 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n79 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n138 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U74  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n12 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n3 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n13 ), .C2(n17297), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n14 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N145 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U75  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n6 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n15 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n8 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n16 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n10 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n17 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n14 ) );
  NOR2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U37  ( .A1(n17112), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n95 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N153 ) );
  NOR2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U38  ( .A1(n17112), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n80 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N154 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U166  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n30 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n38 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n80 ), .C2(n17297), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n81 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N138 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U167  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n10 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n7 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n41 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n82 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n8 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n33 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n81 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U168  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n44 ), .B2(n17102), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n21 ), .C2(n17077), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n87 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n82 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U169  ( .A1(n12649), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n26 ), .B1(
        \pipeline/stageE/input1_to_ALU [1]), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n27 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n87 ) );
  AOI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U106  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n11 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n73 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n9 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n72 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n93 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n80 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U108  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n92 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n67 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n76 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n71 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n94 ) );
  NOR2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U33  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n25 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N159 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U162  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n18 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n38 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n39 ), .C2(n17297), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n40 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N140 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U163  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n10 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n22 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n41 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n42 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n8 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n21 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n40 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U164  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n44 ), .B2(n17088), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n21 ), .C2(n17087), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n48 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n42 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U165  ( .A1(
        \pipeline/stageE/input1_to_ALU [4]), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n26 ), .B1(
        \pipeline/stageE/input1_to_ALU [3]), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n27 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n48 ) );
  AOI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U178  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n51 ), .B2(
        \pipeline/stageE/input1_to_ALU [10]), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n167 ), .C2(
        \pipeline/stageE/input1_to_ALU [9]), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n53 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n18 ) );
  OAI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U179  ( .A1(n17095), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n55 ), .B1(n17089), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n57 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n53 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U158  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n24 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n38 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n60 ), .C2(n17297), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n61 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N139 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U159  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n10 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n28 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n41 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n62 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n8 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n27 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n61 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U160  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n44 ), .B2(n17087), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n21 ), .C2(n17102), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n65 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n62 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U161  ( .A1(
        \pipeline/stageE/input1_to_ALU [3]), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n26 ), .B1(n12649), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n50 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n65 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U72  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n24 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n3 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n25 ), .C2(n17297), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n26 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N143 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U73  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n6 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n27 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n8 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n28 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n10 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n29 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n26 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U127  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n44 ), .B2(n17079), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n21 ), .C2(n17738), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n142 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n28 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U128  ( .A1(
        \pipeline/stageE/input1_to_ALU [15]), .A2(n17110), .B1(
        \pipeline/stageE/input1_to_ALU [14]), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n50 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n142 ) );
  OAI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U148  ( .A1(n17082), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n55 ), .B1(n17085), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n57 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n144 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U55  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n78 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n73 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n59 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n76 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n79 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n72 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n25 ) );
  AOI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U176  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n51 ), .B2(
        \pipeline/stageE/input1_to_ALU [9]), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n167 ), .C2(
        \pipeline/stageE/input1_to_ALU [8]), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n66 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n24 ) );
  OAI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U177  ( .A1(n17089), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n55 ), .B1(n17088), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n57 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n66 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U66  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n30 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n3 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n31 ), .C2(n17297), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n32 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N142 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U67  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n6 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n33 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n8 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n7 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n10 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n9 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n32 ) );
  AOI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U149  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n51 ), .B2(
        \pipeline/stageE/input1_to_ALU [12]), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n167 ), .C2(
        \pipeline/stageE/input1_to_ALU [11]), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n83 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n2 ) );
  OAI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U150  ( .A1(n17085), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n55 ), .B1(n17090), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n57 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n83 ) );
  AOI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U180  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n51 ), .B2(
        \pipeline/stageE/input1_to_ALU [8]), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n167 ), .C2(
        \pipeline/stageE/input1_to_ALU [7]), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n88 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n30 ) );
  OAI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U181  ( .A1(n17088), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n55 ), .B1(n17087), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n57 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n88 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U68  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n34 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n3 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n35 ), .C2(n17297), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n36 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N141 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U69  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n6 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n37 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n8 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n15 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n10 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n16 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n36 ) );
  NOR2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U40  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n13 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N161 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U92  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n74 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n72 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n68 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n73 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n13 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U83  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n96 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n38 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n97 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n3 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n98 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N152 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U85  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n10 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n75 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n99 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n58 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n8 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n77 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n98 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U79  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n103 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n38 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n104 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n3 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n105 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N150 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U82  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n10 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n71 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n99 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n67 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n8 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n11 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n105 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U125  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n44 ), .B2(n17738), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n46 ), .C2(n17101), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n117 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n7 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U126  ( .A1(
        \pipeline/stageE/input1_to_ALU [14]), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n26 ), .B1(n17160), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n50 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n117 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U119  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n44 ), .B2(n17118), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n21 ), .C2(n17097), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n120 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n9 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U120  ( .A1(
        \pipeline/stageE/input1_to_ALU [18]), .A2(n17110), .B1(
        \pipeline/stageE/input1_to_ALU [17]), .B2(n17111), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n120 ) );
  NOR2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U39  ( .A1(n17112), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n60 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N155 ) );
  AOI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U109  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n79 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n73 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n29 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n72 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n90 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n60 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U111  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n92 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n59 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n76 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n78 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n91 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U121  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n44 ), .B2(n17084), .C1(n17118), 
        .C2(\pipeline/stageE/EXE_ALU/alu_shift/C50/n46 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n141 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n29 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U122  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n49 ), .A2(
        \pipeline/stageE/input1_to_ALU [19]), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n50 ), .B2(
        \pipeline/stageE/input1_to_ALU [18]), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n141 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U141  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n44 ), .B2(n17115), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n21 ), .C2(n17117), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n139 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n79 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U142  ( .A1(
        \pipeline/stageE/input1_to_ALU [23]), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n49 ), .B1(
        \pipeline/stageE/input1_to_ALU [22]), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n50 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n139 ) );
  AOI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U103  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n16 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n6 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n15 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n41 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n122 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n121 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U105  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n10 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n74 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n99 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n68 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n8 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n17 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n123 ) );
  NOR2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U13  ( .A1(n17297), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n124 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n99 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U76  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n97 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n38 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n43 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n3 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n125 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N148 ) );
  AOI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U77  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n10 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n77 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n8 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n23 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n126 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n125 ) );
  NOR3_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U78  ( .A1(n17297), .A2(
        n17296), .A3(\pipeline/stageE/EXE_ALU/alu_shift/C50/n69 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n126 ) );
  OAI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U154  ( .A1(n17080), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n55 ), .B1(n17082), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n57 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n132 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U151  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n44 ), .B2(n17096), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n21 ), .C2(n17079), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n137 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n22 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U152  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/A[16] ), .A2(n17110), .B1(
        \pipeline/stageE/input1_to_ALU [15]), .B2(n17111), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n137 ) );
  NOR2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U32  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n31 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N158 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U54  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n71 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n73 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n67 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n76 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n11 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n72 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n31 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U138  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n44 ), .B2(n17117), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n46 ), .C2(n17092), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n108 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n11 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U140  ( .A1(
        \pipeline/stageE/input1_to_ALU [22]), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n49 ), .B1(
        \pipeline/stageE/input1_to_ALU [21]), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n50 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n108 ) );
  NOR2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U31  ( .A1(n17112), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n35 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N157 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U53  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n74 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n73 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n68 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n76 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n17 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n72 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n35 ) );
  NOR2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U36  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n39 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N156 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U57  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n23 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n72 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n77 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n73 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n89 ), .C2(n17296), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n39 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U117  ( .B1(n17118), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n55 ), .C1(n17097), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n57 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n128 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n23 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U118  ( .A1(
        \pipeline/stageE/input1_to_ALU [22]), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n51 ), .B1(
        \pipeline/stageE/input1_to_ALU [21]), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n167 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n128 ) );
  NOR2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U35  ( .A1(n17112), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n4 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N162 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U90  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n71 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n72 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n67 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n73 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n4 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U132  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n44 ), .B2(n17093), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n46 ), .C2(n17078), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n114 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n71 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U133  ( .A1(
        \pipeline/stageE/input1_to_ALU [26]), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n49 ), .B1(
        \pipeline/stageE/input1_to_ALU [25]), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n50 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n114 ) );
  NOR2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U34  ( .A1(n17112), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n19 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N160 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U56  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n75 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n73 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n58 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n76 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n77 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n72 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n19 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U145  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n44 ), .B2(n17086), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n46 ), .C2(n17115), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n131 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n77 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U146  ( .A1(
        \pipeline/stageE/input1_to_ALU [24]), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n49 ), .B1(
        \pipeline/stageE/input1_to_ALU [23]), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n50 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n131 ) );
  NOR2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U41  ( .A1(n17112), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n70 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N163 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U91  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n78 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n72 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n59 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n73 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n70 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U134  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n44 ), .B2(n17094), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n46 ), .C2(n17093), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n143 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n78 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U135  ( .A1(
        \pipeline/stageE/input1_to_ALU [27]), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n49 ), .B1(
        \pipeline/stageE/input1_to_ALU [26]), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n50 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n143 ) );
  NOR3_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U15  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n69 ), .A2(n17112), .A3(n17296), 
        .ZN(\pipeline/stageE/EXE_ALU/alu_shift/N164 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U156  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n44 ), .B2(n17083), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n21 ), .C2(n17094), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n127 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n75 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U157  ( .A1(
        \pipeline/stageE/input1_to_ALU [28]), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n49 ), .B1(
        \pipeline/stageE/input1_to_ALU [27]), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n27 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n127 ) );
  OAI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U51  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n55 ), .A2(n17083), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n46 ), .B2(n17104), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n57 ), .C2(n17094), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n67 ) );
  OAI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U52  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n57 ), .A2(n17083), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n55 ), .B2(n17104), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n59 ) );
  NOR2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U93  ( .A1(n17104), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n57 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n58 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U170  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n34 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n38 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n95 ), .C2(n17297), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n145 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N137 ) );
  AOI222_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U171  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n10 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n15 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n41 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n146 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n8 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n37 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n145 ) );
  AOI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U174  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n51 ), .B2(
        \pipeline/stageE/input1_to_ALU [11]), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n167 ), .C2(
        \pipeline/stageE/input1_to_ALU [10]), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n147 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n12 ) );
  OAI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U175  ( .A1(n17090), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n55 ), .B1(n17095), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n57 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n147 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U172  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n44 ), .B2(n17077), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n46 ), .C2(n17091), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n151 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n146 ) );
  NAND2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U6  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n72 ), .A2(n17297), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n3 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U129  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n44 ), .B2(n17101), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n46 ), .C2(n17100), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n153 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n15 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U131  ( .A1(n17160), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n49 ), .B1(
        \pipeline/stageE/input1_to_ALU [12]), .B2(n17111), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n153 ) );
  NOR2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U28  ( .A1(n17739), .A2(
        n17112), .ZN(\pipeline/stageE/EXE_ALU/alu_shift/C50/n148 ) );
  AOI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U58  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n17 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n73 ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n16 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n72 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n155 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n95 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U60  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n92 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n68 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n76 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n74 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n156 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U136  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n44 ), .B2(n17078), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n46 ), .C2(n17086), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n157 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n74 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U137  ( .A1(
        \pipeline/stageE/input1_to_ALU [25]), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n49 ), .B1(
        \pipeline/stageE/input1_to_ALU [24]), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n50 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n157 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U115  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n44 ), .B2(n17104), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n21 ), .C2(n17083), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n158 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n68 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U116  ( .A1(
        \pipeline/stageE/input1_to_ALU [29]), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n49 ), .B1(
        \pipeline/stageE/input1_to_ALU [28]), .B2(n17111), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n158 ) );
  NOR2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U23  ( .A1(n17081), .A2(
        n17739), .ZN(\pipeline/stageE/EXE_ALU/alu_shift/C50/n92 ) );
  NAND2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U27  ( .A1(n17081), .A2(
        n17739), .ZN(\pipeline/stageE/EXE_ALU/alu_shift/C50/n124 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U123  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n44 ), .B2(n17097), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n21 ), .C2(n17096), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n159 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n16 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U124  ( .A1(
        \pipeline/stageE/input1_to_ALU [17]), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n49 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/A[16] ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n50 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n159 ) );
  OAI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U143  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n55 ), .B2(n17084), .C1(n17118), 
        .C2(\pipeline/stageE/EXE_ALU/alu_shift/C50/n57 ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n160 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n17 ) );
  AOI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U144  ( .A1(
        \pipeline/stageE/input1_to_ALU [23]), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n51 ), .B1(
        \pipeline/stageE/input1_to_ALU [22]), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n167 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n160 ) );
  NAND2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U12  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n73 ), .A2(n17297), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n38 ) );
  AOI221_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U182  ( .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n51 ), .B2(
        \pipeline/stageE/input1_to_ALU [7]), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n167 ), .C2(
        \pipeline/stageE/input1_to_ALU [6]), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n161 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n34 ) );
  OAI22_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U183  ( .A1(n17087), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n55 ), .B1(n17102), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n57 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n161 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C50/U102  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n75 ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n58 ), .S(n17074), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n89 ) );
  AND2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/U38  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][14] ), .A2(n17737), 
        .ZN(\pipeline/stageE/EXE_ALU/alu_shift/N248 ) );
  AND2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/U33  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][9] ), .A2(n17297), 
        .ZN(\pipeline/stageE/EXE_ALU/alu_shift/N243 ) );
  AND2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/U35  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][10] ), .A2(n17302), 
        .ZN(\pipeline/stageE/EXE_ALU/alu_shift/N244 ) );
  AND2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/U39  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][8] ), .A2(n17302), 
        .ZN(\pipeline/stageE/EXE_ALU/alu_shift/N242 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/U13  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/n10 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][0] ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/U10  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/n9 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][1] ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/U16  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/n4 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][6] ) );
  AND2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/U37  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][15] ), .A2(n17302), 
        .ZN(\pipeline/stageE/EXE_ALU/alu_shift/N249 ) );
  AND2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/U36  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][13] ), .A2(n17297), 
        .ZN(\pipeline/stageE/EXE_ALU/alu_shift/N247 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/U11  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/n8 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][2] ) );
  AND2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/U32  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][12] ), .A2(n17302), 
        .ZN(\pipeline/stageE/EXE_ALU/alu_shift/N246 ) );
  AND2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/U34  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][11] ), .A2(n17297), 
        .ZN(\pipeline/stageE/EXE_ALU/alu_shift/N245 ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/U15  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/n5 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][5] ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/U14  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/n6 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][4] ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/U12  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/n7 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][3] ) );
  AND2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/U29  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][1] ), .A2(n17081), 
        .ZN(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][1] ) );
  INV_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/U17  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/n3 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][7] ) );
  AND2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/U30  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][2] ), .A2(n17081), 
        .ZN(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][2] ) );
  AND2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/U31  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][3] ), .A2(n17081), 
        .ZN(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][3] ) );
  AND2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/U46  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][1] ), .A2(n17303), 
        .ZN(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][1] ) );
  AND2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/U44  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][0] ), .A2(n17081), 
        .ZN(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][0] ) );
  AND2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/U48  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][0] ), .A2(n17303), 
        .ZN(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][0] ) );
  NOR2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/U6  ( .A1(n17112), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/n3 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N241 ) );
  NOR2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/U18  ( .A1(n17112), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/n9 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N235 ) );
  NAND2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/U28  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][1] ), .A2(n17739), 
        .ZN(\pipeline/stageE/EXE_ALU/alu_shift/C88/n9 ) );
  NOR2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/U9  ( .A1(n17112), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/n7 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N237 ) );
  NOR2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/U8  ( .A1(n17112), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/n8 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N236 ) );
  NOR2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/U7  ( .A1(n17112), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/n4 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N240 ) );
  NAND2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/U25  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][6] ), .A2(n17739), 
        .ZN(\pipeline/stageE/EXE_ALU/alu_shift/C88/n4 ) );
  NOR2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/U4  ( .A1(n17112), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/n5 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N239 ) );
  NOR2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/U5  ( .A1(n17112), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/n6 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N238 ) );
  NAND2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/U26  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][2] ), .A2(n17739), 
        .ZN(\pipeline/stageE/EXE_ALU/alu_shift/C88/n8 ) );
  NAND2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/U22  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][5] ), .A2(n17739), 
        .ZN(\pipeline/stageE/EXE_ALU/alu_shift/C88/n5 ) );
  NAND2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/U23  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][4] ), .A2(n17739), 
        .ZN(\pipeline/stageE/EXE_ALU/alu_shift/C88/n6 ) );
  NAND2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/U27  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][3] ), .A2(n17739), 
        .ZN(\pipeline/stageE/EXE_ALU/alu_shift/C88/n7 ) );
  NAND2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/U24  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][7] ), .A2(n17739), 
        .ZN(\pipeline/stageE/EXE_ALU/alu_shift/C88/n3 ) );
  NOR2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/U19  ( .A1(n17112), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/n10 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N234 ) );
  NAND2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/U43  ( .A1(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][0] ), .A2(n17739), 
        .ZN(\pipeline/stageE/EXE_ALU/alu_shift/C88/n10 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_0_1  ( .A(
        \pipeline/stageE/input1_to_ALU [1]), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/N202 ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][1] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_0_2  ( .A(n12649), .B(
        \pipeline/stageE/input1_to_ALU [1]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][2] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_0_3  ( .A(
        \pipeline/stageE/input1_to_ALU [3]), .B(n12649), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][3] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_0_4  ( .A(
        \pipeline/stageE/input1_to_ALU [4]), .B(
        \pipeline/stageE/input1_to_ALU [3]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][4] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_0_5  ( .A(
        \pipeline/stageE/input1_to_ALU [5]), .B(
        \pipeline/stageE/input1_to_ALU [4]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][5] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_0_6  ( .A(
        \pipeline/stageE/input1_to_ALU [6]), .B(
        \pipeline/stageE/input1_to_ALU [5]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][6] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_0_7  ( .A(
        \pipeline/stageE/input1_to_ALU [7]), .B(
        \pipeline/stageE/input1_to_ALU [6]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][7] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_0_8  ( .A(
        \pipeline/stageE/input1_to_ALU [8]), .B(
        \pipeline/stageE/input1_to_ALU [7]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][8] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_0_9  ( .A(
        \pipeline/stageE/input1_to_ALU [9]), .B(
        \pipeline/stageE/input1_to_ALU [8]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][9] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_0_10  ( .A(
        \pipeline/stageE/input1_to_ALU [10]), .B(
        \pipeline/stageE/input1_to_ALU [9]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][10] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_0_11  ( .A(
        \pipeline/stageE/input1_to_ALU [11]), .B(
        \pipeline/stageE/input1_to_ALU [10]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][11] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_0_12  ( .A(
        \pipeline/stageE/input1_to_ALU [12]), .B(
        \pipeline/stageE/input1_to_ALU [11]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][12] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_0_13  ( .A(
        \pipeline/stageE/input1_to_ALU [13]), .B(
        \pipeline/stageE/input1_to_ALU [12]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][13] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_0_14  ( .A(
        \pipeline/stageE/input1_to_ALU [14]), .B(
        \pipeline/stageE/input1_to_ALU [13]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][14] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_0_15  ( .A(
        \pipeline/stageE/input1_to_ALU [15]), .B(
        \pipeline/stageE/input1_to_ALU [14]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][15] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_0_16  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/A[16] ), .B(
        \pipeline/stageE/input1_to_ALU [15]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][16] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_0_17  ( .A(
        \pipeline/stageE/input1_to_ALU [17]), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/A[16] ), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][17] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_0_18  ( .A(
        \pipeline/stageE/input1_to_ALU [18]), .B(
        \pipeline/stageE/input1_to_ALU [17]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][18] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_0_19  ( .A(
        \pipeline/stageE/input1_to_ALU [19]), .B(
        \pipeline/stageE/input1_to_ALU [18]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][19] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_0_20  ( .A(
        \pipeline/stageE/input1_to_ALU [20]), .B(
        \pipeline/stageE/input1_to_ALU [19]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][20] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_0_21  ( .A(
        \pipeline/stageE/input1_to_ALU [21]), .B(
        \pipeline/stageE/input1_to_ALU [20]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][21] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_0_22  ( .A(
        \pipeline/stageE/input1_to_ALU [22]), .B(
        \pipeline/stageE/input1_to_ALU [21]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][22] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_0_23  ( .A(
        \pipeline/stageE/input1_to_ALU [23]), .B(
        \pipeline/stageE/input1_to_ALU [22]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][23] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_0_24  ( .A(
        \pipeline/stageE/input1_to_ALU [24]), .B(
        \pipeline/stageE/input1_to_ALU [23]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][24] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_0_25  ( .A(
        \pipeline/stageE/input1_to_ALU [25]), .B(
        \pipeline/stageE/input1_to_ALU [24]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][25] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_0_26  ( .A(
        \pipeline/stageE/input1_to_ALU [26]), .B(
        \pipeline/stageE/input1_to_ALU [25]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][26] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_0_27  ( .A(
        \pipeline/stageE/input1_to_ALU [27]), .B(
        \pipeline/stageE/input1_to_ALU [26]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][27] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_0_28  ( .A(
        \pipeline/stageE/input1_to_ALU [28]), .B(
        \pipeline/stageE/input1_to_ALU [27]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][28] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_0_29  ( .A(
        \pipeline/stageE/input1_to_ALU [29]), .B(
        \pipeline/stageE/input1_to_ALU [28]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][29] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_0_30  ( .A(
        \pipeline/stageE/input1_to_ALU [30]), .B(
        \pipeline/stageE/input1_to_ALU [29]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][30] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_0_31  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/N136 ), .B(
        \pipeline/stageE/input1_to_ALU [30]), .S(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][31] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_1_2  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][2] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][0] ), .S(n17099), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][2] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_1_3  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][3] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][1] ), .S(n17099), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][3] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_1_4  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][4] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][2] ), .S(n17099), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][4] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_1_5  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][5] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][3] ), .S(n17099), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][5] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_1_6  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][6] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][4] ), .S(n17099), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][6] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_1_7  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][7] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][5] ), .S(n17099), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][7] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_1_8  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][8] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][6] ), .S(n17099), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][8] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_1_9  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][9] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][7] ), .S(n17099), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][9] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_1_10  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][10] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][8] ), .S(n17099), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][10] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_1_11  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][11] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][9] ), .S(n17099), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][11] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_1_12  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][12] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][10] ), .S(n17099), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][12] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_1_13  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][13] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][11] ), .S(n17099), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][13] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_1_14  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][14] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][12] ), .S(n17099), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][14] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_1_15  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][15] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][13] ), .S(n17099), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][15] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_1_16  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][16] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][14] ), .S(n17099), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][16] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_1_17  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][17] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][15] ), .S(n17099), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][17] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_1_18  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][18] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][16] ), .S(n17099), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][18] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_1_19  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][19] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][17] ), .S(n17099), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][19] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_1_20  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][20] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][18] ), .S(n17099), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][20] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_1_21  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][21] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][19] ), .S(n17099), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][21] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_1_22  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][22] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][20] ), .S(n17099), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][22] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_1_23  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][23] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][21] ), .S(n17099), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][23] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_1_24  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][24] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][22] ), .S(n17099), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][24] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_1_25  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][25] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][23] ), .S(n17099), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][25] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_1_26  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][26] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][24] ), .S(n17099), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][26] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_1_27  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][27] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][25] ), .S(n17099), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][27] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_1_28  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][28] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][26] ), .S(n17099), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][28] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_1_29  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][29] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][27] ), .S(n17099), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][29] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_1_30  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][30] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][28] ), .S(n17099), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][30] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_1_31  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][31] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][29] ), .S(n17099), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][31] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_2_4  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][4] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][0] ), .S(n17114), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][4] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_2_5  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][5] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][1] ), .S(n17114), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][5] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_2_6  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][6] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][2] ), .S(n17114), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][6] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_2_7  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][7] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][3] ), .S(n17114), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][7] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_2_8  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][8] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][4] ), .S(n17114), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][8] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_2_9  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][9] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][5] ), .S(n17114), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][9] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_2_10  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][10] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][6] ), .S(n17114), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][10] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_2_11  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][11] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][7] ), .S(n17114), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][11] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_2_12  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][12] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][8] ), .S(n17114), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][12] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_2_13  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][13] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][9] ), .S(n17114), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][13] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_2_14  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][14] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][10] ), .S(n17114), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][14] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_2_15  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][15] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][11] ), .S(n17114), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][15] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_2_16  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][16] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][12] ), .S(n17114), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][16] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_2_17  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][17] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][13] ), .S(n17114), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][17] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_2_18  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][18] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][14] ), .S(n17114), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][18] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_2_19  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][19] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][15] ), .S(n17114), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][19] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_2_20  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][20] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][16] ), .S(n17114), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][20] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_2_21  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][21] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][17] ), .S(n17114), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][21] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_2_22  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][22] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][18] ), .S(n17114), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][22] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_2_23  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][23] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][19] ), .S(n17114), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][23] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_2_24  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][24] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][20] ), .S(n17114), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][24] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_2_25  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][25] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][21] ), .S(n17114), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][25] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_2_26  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][26] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][22] ), .S(n17114), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][26] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_2_27  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][27] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][23] ), .S(n17114), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][27] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_2_28  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][28] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][24] ), .S(n17114), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][28] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_2_29  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][29] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][25] ), .S(n17114), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][29] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_2_30  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][30] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][26] ), .S(n17114), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][30] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_2_31  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][31] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[2][27] ), .S(n17114), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][31] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_3_8  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][8] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][0] ), .S(n17296), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][8] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_3_9  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][9] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][1] ), .S(n17301), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][9] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_3_10  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][10] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][2] ), .S(n17300), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][10] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_3_11  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][11] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][3] ), .S(n17301), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][11] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_3_12  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][12] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][4] ), .S(n17301), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][12] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_3_13  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][13] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][5] ), .S(n17300), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][13] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_3_14  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][14] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][6] ), .S(n17300), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][14] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_3_15  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][15] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][7] ), .S(n17299), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][15] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_3_16  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][16] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][8] ), .S(n17296), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][16] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_3_17  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][17] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][9] ), .S(n17299), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][17] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_3_18  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][18] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][10] ), .S(n17301), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][18] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_3_19  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][19] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][11] ), .S(n17296), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][19] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_3_20  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][20] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][12] ), .S(n17300), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][20] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_3_21  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][21] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][13] ), .S(n17296), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][21] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_3_22  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][22] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][14] ), .S(n17300), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][22] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_3_23  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][23] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][15] ), .S(n17301), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][23] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_3_24  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][24] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][16] ), .S(n17301), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][24] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_3_25  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][25] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][17] ), .S(n17299), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][25] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_3_26  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][26] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][18] ), .S(n17300), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][26] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_3_27  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][27] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][19] ), .S(n17296), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][27] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_3_28  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][28] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][20] ), .S(n17300), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][28] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_3_29  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][29] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][21] ), .S(n17301), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][29] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_3_30  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][30] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][22] ), .S(n17299), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][30] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_3_31  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][31] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[3][23] ), .S(n17299), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][31] ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_4_16  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][16] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][0] ), .S(n17112), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N250 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_4_17  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][17] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][1] ), .S(n17112), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N251 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_4_18  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][18] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][2] ), .S(n17112), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N252 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_4_19  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][19] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][3] ), .S(n17112), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N253 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_4_20  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][20] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][4] ), .S(n17112), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N254 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_4_21  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][21] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][5] ), .S(n17112), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N255 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_4_22  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][22] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][6] ), .S(n17112), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N256 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_4_23  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][23] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][7] ), .S(n17112), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N257 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_4_24  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][24] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][8] ), .S(n17112), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N258 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_4_25  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][25] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][9] ), .S(n17112), .Z(
        \pipeline/stageE/EXE_ALU/alu_shift/N259 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_4_26  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][26] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][10] ), .S(n17112), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/N260 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_4_27  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][27] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][11] ), .S(n17112), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/N261 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_4_28  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][28] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][12] ), .S(n17112), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/N262 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_4_29  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][29] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][13] ), .S(n17112), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/N263 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_4_30  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][30] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][14] ), .S(n17112), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/N264 ) );
  MUX2_X1 \pipeline/stageE/EXE_ALU/alu_shift/C88/M1_4_31  ( .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][31] ), .B(
        \pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[4][15] ), .S(n17112), 
        .Z(\pipeline/stageE/EXE_ALU/alu_shift/N265 ) );
  INV_X1 \pipeline/stageD/evaluate_jump_target/add_29/U41  ( .A(
        \pipeline/stageD/offset_to_jump_temp [24]), .ZN(
        \pipeline/stageD/evaluate_jump_target/add_29/n168 ) );
  INV_X1 \pipeline/stageD/evaluate_jump_target/add_29/U57  ( .A(
        \pipeline/stageD/offset_to_jump_temp [20]), .ZN(
        \pipeline/stageD/evaluate_jump_target/add_29/n180 ) );
  INV_X1 \pipeline/stageD/evaluate_jump_target/add_29/U75  ( .A(
        \pipeline/stageD/offset_to_jump_temp [16]), .ZN(
        \pipeline/stageD/evaluate_jump_target/add_29/n194 ) );
  INV_X1 \pipeline/stageD/evaluate_jump_target/add_29/U67  ( .A(
        \pipeline/stageD/offset_to_jump_temp [18]), .ZN(
        \pipeline/stageD/evaluate_jump_target/add_29/n188 ) );
  INV_X1 \pipeline/stageD/evaluate_jump_target/add_29/U49  ( .A(
        \pipeline/stageD/offset_to_jump_temp [22]), .ZN(
        \pipeline/stageD/evaluate_jump_target/add_29/n174 ) );
  XNOR2_X1 \pipeline/stageD/evaluate_jump_target/add_29/U59  ( .A(
        \pipeline/stageD/evaluate_jump_target/add_29/n183 ), .B(
        \pipeline/stageD/evaluate_jump_target/add_29/n184 ), .ZN(
        \pipeline/stageD/evaluate_jump_target/N34 ) );
  XNOR2_X1 \pipeline/stageD/evaluate_jump_target/add_29/U14  ( .A(
        \pipeline/nextPC_IFID_DEC[3] ), .B(
        \pipeline/stageD/offset_to_jump_temp [3]), .ZN(
        \pipeline/stageD/evaluate_jump_target/add_29/n144 ) );
  XNOR2_X1 \pipeline/stageD/evaluate_jump_target/add_29/U10  ( .A(
        \pipeline/nextPC_IFID_DEC[5] ), .B(
        \pipeline/stageD/offset_to_jump_temp [5]), .ZN(
        \pipeline/stageD/evaluate_jump_target/add_29/n138 ) );
  AOI22_X1 \pipeline/stageD/evaluate_jump_target/add_29/U12  ( .A1(
        \pipeline/nextPC_IFID_DEC[4] ), .A2(
        \pipeline/stageD/offset_to_jump_temp [4]), .B1(n17412), .B2(n17455), 
        .ZN(\pipeline/stageD/evaluate_jump_target/add_29/n141 ) );
  AOI22_X1 \pipeline/stageD/evaluate_jump_target/add_29/U8  ( .A1(
        \pipeline/nextPC_IFID_DEC[6] ), .A2(
        \pipeline/stageD/offset_to_jump_temp [6]), .B1(n17361), .B2(n17456), 
        .ZN(\pipeline/stageD/evaluate_jump_target/add_29/n135 ) );
  XNOR2_X1 \pipeline/stageD/evaluate_jump_target/add_29/U6  ( .A(
        \pipeline/nextPC_IFID_DEC[7] ), .B(
        \pipeline/stageD/offset_to_jump_temp [7]), .ZN(
        \pipeline/stageD/evaluate_jump_target/add_29/n132 ) );
  AOI22_X1 \pipeline/stageD/evaluate_jump_target/add_29/U4  ( .A1(
        \pipeline/nextPC_IFID_DEC[8] ), .A2(
        \pipeline/stageD/offset_to_jump_temp [8]), .B1(n17428), .B2(n17457), 
        .ZN(\pipeline/stageD/evaluate_jump_target/add_29/n129 ) );
  XNOR2_X1 \pipeline/stageD/evaluate_jump_target/add_29/U2  ( .A(
        \pipeline/stageD/offset_to_jump_temp [9]), .B(
        \pipeline/nextPC_IFID_DEC[9] ), .ZN(
        \pipeline/stageD/evaluate_jump_target/add_29/n126 ) );
  AOI22_X1 \pipeline/stageD/evaluate_jump_target/add_29/U97  ( .A1(
        \pipeline/nextPC_IFID_DEC[10] ), .A2(
        \pipeline/stageD/offset_to_jump_temp [10]), .B1(n17440), .B2(n17458), 
        .ZN(\pipeline/stageD/evaluate_jump_target/add_29/n213 ) );
  XNOR2_X1 \pipeline/stageD/evaluate_jump_target/add_29/U93  ( .A(
        \pipeline/stageD/evaluate_jump_target/add_29/n209 ), .B(n17174), .ZN(
        \pipeline/stageD/evaluate_jump_target/N44 ) );
  XNOR2_X1 \pipeline/stageD/evaluate_jump_target/add_29/U95  ( .A(
        \pipeline/nextPC_IFID_DEC[11] ), .B(
        \pipeline/stageD/offset_to_jump_temp [11]), .ZN(
        \pipeline/stageD/evaluate_jump_target/add_29/n209 ) );
  XNOR2_X1 \pipeline/stageD/evaluate_jump_target/add_29/U88  ( .A(n17178), .B(
        \pipeline/stageD/evaluate_jump_target/add_29/n207 ), .ZN(
        \pipeline/stageD/evaluate_jump_target/N45 ) );
  AOI22_X1 \pipeline/stageD/evaluate_jump_target/add_29/U89  ( .A1(
        \pipeline/nextPC_IFID_DEC[12] ), .A2(
        \pipeline/stageD/offset_to_jump_temp [12]), .B1(n17444), .B2(n17459), 
        .ZN(\pipeline/stageD/evaluate_jump_target/add_29/n207 ) );
  XNOR2_X1 \pipeline/stageD/evaluate_jump_target/add_29/U87  ( .A(
        \pipeline/nextPC_IFID_DEC[13] ), .B(
        \pipeline/stageD/offset_to_jump_temp [13]), .ZN(
        \pipeline/stageD/evaluate_jump_target/add_29/n203 ) );
  AOI22_X1 \pipeline/stageD/evaluate_jump_target/add_29/U81  ( .A1(
        \pipeline/nextPC_IFID_DEC[14] ), .A2(
        \pipeline/stageD/offset_to_jump_temp [14]), .B1(n17445), .B2(n17460), 
        .ZN(\pipeline/stageD/evaluate_jump_target/add_29/n201 ) );
  XNOR2_X1 \pipeline/stageD/evaluate_jump_target/add_29/U79  ( .A(
        \pipeline/nextPC_IFID_DEC[15] ), .B(
        \pipeline/stageD/offset_to_jump_temp [15]), .ZN(
        \pipeline/stageD/evaluate_jump_target/add_29/n197 ) );
  AOI22_X1 \pipeline/stageD/evaluate_jump_target/add_29/U73  ( .A1(
        \pipeline/nextPC_IFID_DEC[16] ), .A2(
        \pipeline/stageD/offset_to_jump_temp [16]), .B1(
        \pipeline/stageD/evaluate_jump_target/add_29/n194 ), .B2(n17461), .ZN(
        \pipeline/stageD/evaluate_jump_target/add_29/n195 ) );
  XNOR2_X1 \pipeline/stageD/evaluate_jump_target/add_29/U71  ( .A(
        \pipeline/nextPC_IFID_DEC[17] ), .B(
        \pipeline/stageD/offset_to_jump_temp [17]), .ZN(
        \pipeline/stageD/evaluate_jump_target/add_29/n191 ) );
  AOI22_X1 \pipeline/stageD/evaluate_jump_target/add_29/U65  ( .A1(
        \pipeline/nextPC_IFID_DEC[18] ), .A2(
        \pipeline/stageD/offset_to_jump_temp [18]), .B1(
        \pipeline/stageD/evaluate_jump_target/add_29/n188 ), .B2(n17462), .ZN(
        \pipeline/stageD/evaluate_jump_target/add_29/n189 ) );
  XNOR2_X1 \pipeline/stageD/evaluate_jump_target/add_29/U63  ( .A(
        \pipeline/nextPC_IFID_DEC[19] ), .B(
        \pipeline/stageD/offset_to_jump_temp [19]), .ZN(
        \pipeline/stageD/evaluate_jump_target/add_29/n185 ) );
  AOI22_X1 \pipeline/stageD/evaluate_jump_target/add_29/U55  ( .A1(
        \pipeline/nextPC_IFID_DEC[20] ), .A2(
        \pipeline/stageD/offset_to_jump_temp [20]), .B1(
        \pipeline/stageD/evaluate_jump_target/add_29/n180 ), .B2(n17463), .ZN(
        \pipeline/stageD/evaluate_jump_target/add_29/n181 ) );
  XNOR2_X1 \pipeline/stageD/evaluate_jump_target/add_29/U53  ( .A(
        \pipeline/nextPC_IFID_DEC[21] ), .B(
        \pipeline/stageD/offset_to_jump_temp [21]), .ZN(
        \pipeline/stageD/evaluate_jump_target/add_29/n177 ) );
  AOI22_X1 \pipeline/stageD/evaluate_jump_target/add_29/U47  ( .A1(
        \pipeline/nextPC_IFID_DEC[22] ), .A2(
        \pipeline/stageD/offset_to_jump_temp [22]), .B1(
        \pipeline/stageD/evaluate_jump_target/add_29/n174 ), .B2(n17464), .ZN(
        \pipeline/stageD/evaluate_jump_target/add_29/n175 ) );
  XNOR2_X1 \pipeline/stageD/evaluate_jump_target/add_29/U45  ( .A(
        \pipeline/nextPC_IFID_DEC[23] ), .B(
        \pipeline/stageD/offset_to_jump_temp [23]), .ZN(
        \pipeline/stageD/evaluate_jump_target/add_29/n171 ) );
  AOI22_X1 \pipeline/stageD/evaluate_jump_target/add_29/U39  ( .A1(
        \pipeline/nextPC_IFID_DEC[24] ), .A2(
        \pipeline/stageD/offset_to_jump_temp [24]), .B1(
        \pipeline/stageD/evaluate_jump_target/add_29/n168 ), .B2(n17465), .ZN(
        \pipeline/stageD/evaluate_jump_target/add_29/n169 ) );
  XNOR2_X1 \pipeline/stageD/evaluate_jump_target/add_29/U37  ( .A(
        \pipeline/nextPC_IFID_DEC[25] ), .B(
        \pipeline/stageD/offset_to_jump_temp [30]), .ZN(
        \pipeline/stageD/evaluate_jump_target/add_29/n165 ) );
  AOI22_X1 \pipeline/stageD/evaluate_jump_target/add_29/U31  ( .A1(
        \pipeline/nextPC_IFID_DEC[26] ), .A2(
        \pipeline/stageD/offset_to_jump_temp [30]), .B1(n17200), .B2(n17466), 
        .ZN(\pipeline/stageD/evaluate_jump_target/add_29/n163 ) );
  XNOR2_X1 \pipeline/stageD/evaluate_jump_target/add_29/U29  ( .A(
        \pipeline/nextPC_IFID_DEC[27] ), .B(
        \pipeline/stageD/offset_to_jump_temp [30]), .ZN(
        \pipeline/stageD/evaluate_jump_target/add_29/n159 ) );
  AOI22_X1 \pipeline/stageD/evaluate_jump_target/add_29/U23  ( .A1(
        \pipeline/nextPC_IFID_DEC[28] ), .A2(
        \pipeline/stageD/offset_to_jump_temp [30]), .B1(n17200), .B2(n17467), 
        .ZN(\pipeline/stageD/evaluate_jump_target/add_29/n157 ) );
  XOR2_X1 \pipeline/stageD/evaluate_jump_target/add_29/U120  ( .A(net175543), 
        .B(\pipeline/nextPC_IFID_DEC[0] ), .Z(
        \pipeline/stageD/evaluate_jump_target/N33 ) );
  XOR2_X1 \pipeline/stageD/evaluate_jump_target/add_29/U119  ( .A(
        \pipeline/nextPC_IFID_DEC[1] ), .B(
        \pipeline/stageD/offset_to_jump_temp [1]), .Z(
        \pipeline/stageD/evaluate_jump_target/add_29/n184 ) );
  NOR2_X1 U10950 ( .A1(\pipeline/inst_IFID_DEC[31] ), .A2(
        \pipeline/inst_IFID_DEC[28] ), .ZN(n14190) );
  NAND2_X1 U10948 ( .A1(n14190), .A2(n17382), .ZN(n14177) );
  NOR3_X1 U10947 ( .A1(n13281), .A2(n17313), .A3(n14177), .ZN(n13979) );
  INV_X1 U11908 ( .A(addr_to_dataRam[2]), .ZN(n17012) );
  NAND2_X1 U11734 ( .A1(addr_to_dataRam[4]), .A2(addr_to_dataRam[3]), .ZN(
        n17013) );
  INV_X1 U11873 ( .A(addr_to_dataRam[3]), .ZN(n17015) );
  OAI21_X2 U11253 ( .B1(n17662), .B2(n17321), .A(n16701), .ZN(
        \pipeline/stageE/input1_to_ALU [1]) );
  NOR2_X2 U8598 ( .A1(n13281), .A2(\pipeline/WB_controls_in_MEMWB[0] ), .ZN(
        n14134) );
  NOR2_X2 U9351 ( .A1(n14860), .A2(n14866), .ZN(n14223) );
  NOR2_X2 U9340 ( .A1(n14865), .A2(n14861), .ZN(n14214) );
  NOR2_X2 U9337 ( .A1(n14863), .A2(n14861), .ZN(n14212) );
  NOR2_X2 U9334 ( .A1(n14860), .A2(n14861), .ZN(n14210) );
  NOR2_X2 U9343 ( .A1(n14864), .A2(n14861), .ZN(n14216) );
  NOR3_X1 U10234 ( .A1(n17409), .A2(n17313), .A3(n14177), .ZN(n14947) );
  AND3_X2 U11803 ( .A1(n17012), .A2(n17015), .A3(addr_to_dataRam[4]), .ZN(
        n16822) );
  NAND2_X1 U10243 ( .A1(n17703), .A2(n15646), .ZN(n14168) );
  INV_X1 U10242 ( .A(n14168), .ZN(n14167) );
  DFFR_X1 \pipeline/stageF/PC_reg/PC_out_reg[30]  ( .D(n3989), .CK(Clk), .RN(
        n17703), .Q(n13782), .QN(n7710) );
  DFF_X2 \pipeline/IFID_stage/Instr_out_IFID_reg[1]  ( .D(n3986), .CK(Clk), 
        .Q(\pipeline/stageD/offset_to_jump_temp [1]), .QN(n17406) );
  OAI21_X1 U12262 ( .B1(n14127), .B2(n17018), .A(n17704), .ZN(n14122) );
  OR2_X1 U12263 ( .A1(n14125), .A2(n14126), .ZN(n17018) );
  AOI222_X1 U12264 ( .A1(n15598), .A2(n17579), .B1(n15598), .B2(
        \pipeline/stageE/input1_to_ALU [3]), .C1(n16688), .C2(
        \pipeline/stageE/input1_to_ALU [3]), .ZN(n15566) );
  INV_X1 U12265 ( .A(\pipeline/stageE/input1_to_ALU [30]), .ZN(n17083) );
  INV_X1 U12266 ( .A(\pipeline/stageE/input1_to_ALU [19]), .ZN(n17097) );
  INV_X1 U12267 ( .A(\pipeline/stageE/input1_to_ALU [5]), .ZN(n17087) );
  AND2_X1 U12268 ( .A1(n17019), .A2(n17020), .ZN(n12766) );
  BUF_X2 U12269 ( .A(n12766), .Z(n17155) );
  NOR2_X1 U12270 ( .A1(\pipeline/EXE_controls_in_EXEcute [0]), .A2(n13846), 
        .ZN(n17021) );
  AOI22_X1 U12271 ( .A1(n17666), .A2(\pipeline/Alu_Out_Addr_to_mem[3] ), .B1(
        \pipeline/data_to_RF_from_WB[3] ), .B2(n15123), .ZN(n17022) );
  OAI21_X1 U12272 ( .B1(n17642), .B2(n17021), .A(n17022), .ZN(n17023) );
  OAI21_X2 U12273 ( .B1(\pipeline/immediate_to_exe [3]), .B2(n17327), .A(
        n17023), .ZN(n17739) );
  NAND4_X1 U12274 ( .A1(n15045), .A2(n14970), .A3(n14948), .A4(n15046), .ZN(
        n17024) );
  NOR4_X1 U12275 ( .A1(n15041), .A2(n15042), .A3(n15043), .A4(n17024), .ZN(
        n17025) );
  NAND2_X1 U12276 ( .A1(n17025), .A2(n15037), .ZN(n17026) );
  NOR4_X1 U12277 ( .A1(n15035), .A2(n15033), .A3(n15034), .A4(n17026), .ZN(
        n17027) );
  AND4_X1 U12278 ( .A1(n15039), .A2(n15040), .A3(n17027), .A4(n15032), .ZN(
        n17028) );
  NAND3_X1 U12279 ( .A1(n15030), .A2(n15029), .A3(n17028), .ZN(n17029) );
  NOR4_X1 U12280 ( .A1(n15026), .A2(n15025), .A3(n15027), .A4(n17029), .ZN(
        n17030) );
  NAND2_X1 U12281 ( .A1(n15017), .A2(n17030), .ZN(n17538) );
  AOI21_X1 U12282 ( .B1(n15138), .B2(n15137), .A(n17608), .ZN(n17031) );
  AOI21_X1 U12283 ( .B1(n15142), .B2(n17542), .A(n17031), .ZN(n17032) );
  AOI21_X1 U12284 ( .B1(n17104), .B2(n15137), .A(n17032), .ZN(n15005) );
  OR2_X1 U12285 ( .A1(n17327), .A2(\pipeline/immediate_to_exe [1]), .ZN(n17033) );
  OAI21_X1 U12286 ( .B1(n17642), .B2(n17577), .A(n16699), .ZN(n17034) );
  NAND2_X1 U12287 ( .A1(n17034), .A2(n17033), .ZN(n17741) );
  NOR4_X1 U12288 ( .A1(n15022), .A2(n15021), .A3(n15023), .A4(n15024), .ZN(
        n17035) );
  NAND2_X1 U12289 ( .A1(n15020), .A2(n17035), .ZN(n17537) );
  INV_X1 U12290 ( .A(n17411), .ZN(n17036) );
  NOR3_X1 U12291 ( .A1(\pipeline/EXE_controls_in_EXEcute [2]), .A2(
        \pipeline/EXE_controls_in_EXEcute [4]), .A3(n17036), .ZN(n17528) );
  AOI22_X1 U12292 ( .A1(n17742), .A2(
        \pipeline/stageE/EXE_ALU/add_alu/sCout[0] ), .B1(
        \pipeline/stageE/input2_to_ALU[0] ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/N202 ), .ZN(n15048) );
  AOI22_X1 U12293 ( .A1(n17664), .A2(n13832), .B1(n17663), .B2(
        \pipeline/Alu_Out_Addr_to_mem[5] ), .ZN(n17037) );
  OAI21_X1 U12294 ( .B1(n17105), .B2(n17308), .A(n17037), .ZN(
        \pipeline/stageE/input1_to_ALU [5]) );
  NOR2_X1 U12295 ( .A1(\pipeline/EXE_controls_in_EXEcute [0]), .A2(n13811), 
        .ZN(n17038) );
  OAI21_X1 U12296 ( .B1(n17642), .B2(n17038), .A(n16704), .ZN(n17039) );
  OAI21_X1 U12297 ( .B1(\pipeline/immediate_to_exe [2]), .B2(n17327), .A(
        n17039), .ZN(n17740) );
  OAI21_X1 U12298 ( .B1(n17166), .B2(\pipeline/stageD/offset_to_jump_temp [23]), .A(\pipeline/nextPC_IFID_DEC[23] ), .ZN(n17196) );
  AOI222_X1 U12299 ( .A1(\pipeline/Alu_Out_Addr_to_mem[30] ), .A2(n17331), 
        .B1(n13782), .B2(n17674), .C1(n17108), .C2(
        \pipeline/stageF/PC_plus4/N37 ), .ZN(n17638) );
  AND3_X1 U12300 ( .A1(n15383), .A2(n15368), .A3(n15367), .ZN(n17040) );
  NOR2_X1 U12301 ( .A1(n17040), .A2(n15352), .ZN(n17041) );
  XNOR2_X1 U12302 ( .A(n17041), .B(n17096), .ZN(n17042) );
  XNOR2_X1 U12303 ( .A(n17042), .B(n15348), .ZN(n15021) );
  INV_X1 U12304 ( .A(n17121), .ZN(n17043) );
  AOI222_X1 U12305 ( .A1(n17043), .A2(\pipeline/data_to_RF_from_WB[2] ), .B1(
        n17663), .B2(\pipeline/Alu_Out_Addr_to_mem[2] ), .C1(n16620), .C2(
        n13809), .ZN(n17044) );
  INV_X1 U12306 ( .A(n17044), .ZN(n12649) );
  AOI22_X1 U12307 ( .A1(n17428), .A2(n17457), .B1(
        \pipeline/stageD/evaluate_jump_target/add_29/n128 ), .B2(n17295), .ZN(
        n17177) );
  NOR4_X1 U12308 ( .A1(n16554), .A2(n16796), .A3(n16795), .A4(n17387), .ZN(
        n16619) );
  NAND2_X1 U12309 ( .A1(\pipeline/stageE/input1_to_ALU [23]), .A2(n15263), 
        .ZN(n17045) );
  AOI21_X1 U12310 ( .B1(n15265), .B2(n17045), .A(n17603), .ZN(n17046) );
  NAND2_X1 U12311 ( .A1(n17045), .A2(n15268), .ZN(n17047) );
  OAI21_X1 U12312 ( .B1(n15282), .B2(n17047), .A(n17046), .ZN(n15248) );
  AOI22_X1 U12313 ( .A1(n17739), .A2(n17381), .B1(
        \pipeline/stageE/EXE_ALU/add_alu/sCout[0] ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[3] ), .ZN(n15598) );
  NAND4_X1 U12314 ( .A1(n17279), .A2(n17278), .A3(
        \pipeline/nextPC_IFID_DEC[29] ), .A4(n17183), .ZN(n17186) );
  AOI222_X1 U12315 ( .A1(n15368), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/A[16] ), .B1(n15368), .B2(
        n15369), .C1(\pipeline/stageE/EXE_ALU/alu_shift/C48/A[16] ), .C2(
        n15369), .ZN(n17048) );
  NAND2_X1 U12316 ( .A1(n15367), .A2(n15366), .ZN(n17049) );
  XOR2_X1 U12317 ( .A(n17048), .B(n17049), .Z(n15025) );
  INV_X1 U12318 ( .A(n14094), .ZN(n17050) );
  AOI22_X1 U12319 ( .A1(n14094), .A2(
        \pipeline/stageD/offset_jump_sign_ext [24]), .B1(
        \pipeline/stageD/offset_jump_sign_ext [19]), .B2(n17050), .ZN(n17051)
         );
  AOI22_X1 U12320 ( .A1(n14094), .A2(
        \pipeline/stageD/offset_jump_sign_ext [31]), .B1(
        \pipeline/stageD/offset_jump_sign_ext [20]), .B2(n17050), .ZN(n17052)
         );
  NOR3_X1 U12321 ( .A1(n14091), .A2(n14087), .A3(n14098), .ZN(n17053) );
  OAI22_X1 U12322 ( .A1(n14116), .A2(
        \pipeline/stageD/offset_jump_sign_ext [16]), .B1(
        \pipeline/stageD/offset_jump_sign_ext [17]), .B2(n14117), .ZN(n17054)
         );
  AOI221_X1 U12323 ( .B1(n14116), .B2(
        \pipeline/stageD/offset_jump_sign_ext [16]), .C1(n14117), .C2(
        \pipeline/stageD/offset_jump_sign_ext [17]), .A(n17054), .ZN(n17055)
         );
  OAI211_X1 U12324 ( .C1(n14113), .C2(
        \pipeline/stageD/offset_jump_sign_ext [18]), .A(n17055), .B(n14091), 
        .ZN(n17056) );
  AOI21_X1 U12325 ( .B1(n14113), .B2(
        \pipeline/stageD/offset_jump_sign_ext [18]), .A(n17056), .ZN(n17057)
         );
  XNOR2_X1 U12326 ( .A(n14101), .B(n17052), .ZN(n17058) );
  OAI21_X1 U12327 ( .B1(n17057), .B2(n17053), .A(n17058), .ZN(n17059) );
  XOR2_X1 U12328 ( .A(n14100), .B(n17051), .Z(n17060) );
  NOR3_X1 U12329 ( .A1(n17060), .A2(n14096), .A3(n17059), .ZN(n14092) );
  NAND4_X1 U12330 ( .A1(\pipeline/inst_IFID_DEC[29] ), .A2(n14049), .A3(n13993), .A4(\pipeline/inst_IFID_DEC[27] ), .ZN(n17061) );
  OAI211_X1 U12331 ( .C1(n14059), .C2(n14058), .A(n14020), .B(n17061), .ZN(
        n17062) );
  NOR2_X1 U12332 ( .A1(n17350), .A2(n14064), .ZN(n17063) );
  AOI21_X1 U12333 ( .B1(n14065), .B2(n17076), .A(n17063), .ZN(n17064) );
  AOI221_X1 U12334 ( .B1(n14066), .B2(n17064), .C1(n17076), .C2(n17064), .A(
        n14012), .ZN(n17065) );
  AOI211_X1 U12335 ( .C1(n14032), .C2(n14033), .A(n17062), .B(n17065), .ZN(
        n14041) );
  OAI221_X1 U12336 ( .B1(n15000), .B2(\pipeline/EXE_controls_in_EXEcute [2]), 
        .C1(n15000), .C2(n15001), .A(n17529), .ZN(n17066) );
  AOI21_X1 U12337 ( .B1(n14964), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N105 ), 
        .A(n17623), .ZN(n17067) );
  NAND2_X1 U12338 ( .A1(n17066), .A2(n17067), .ZN(\pipeline/EXMEM_stage/N7 )
         );
  INV_X1 U12339 ( .A(n17106), .ZN(n17068) );
  NAND2_X1 U12340 ( .A1(n17330), .A2(\pipeline/Alu_Out_Addr_to_mem[29] ), .ZN(
        n17069) );
  NAND3_X1 U12341 ( .A1(n17069), .A2(n17622), .A3(n17621), .ZN(n17070) );
  AOI21_X1 U12342 ( .B1(\pipeline/data_to_RF_from_WB[29] ), .B2(n17332), .A(
        n17070), .ZN(n17071) );
  NAND2_X1 U12343 ( .A1(n15607), .A2(\pipeline/stageD/target_Jump_temp [29]), 
        .ZN(n17072) );
  OAI211_X1 U12344 ( .C1(n14887), .C2(n17068), .A(n17071), .B(n17072), .ZN(
        n3988) );
  AND2_X2 U12345 ( .A1(n17233), .A2(n17232), .ZN(n17162) );
  AND2_X2 U12346 ( .A1(n17263), .A2(n17262), .ZN(
        \pipeline/stageD/evaluate_jump_target/add_29/n133 ) );
  INV_X1 U12347 ( .A(n17740), .ZN(n17073) );
  INV_X4 U12348 ( .A(n17740), .ZN(n17074) );
  NOR2_X2 U12349 ( .A1(n16691), .A2(n12649), .ZN(n15055) );
  NAND2_X4 U12350 ( .A1(n14025), .A2(n14167), .ZN(n17075) );
  INV_X2 U12351 ( .A(n4376), .ZN(n17737) );
  NOR2_X4 U12352 ( .A1(n15648), .A2(n15646), .ZN(n15600) );
  BUF_X4 U12353 ( .A(\pipeline/stageE/EXE_ALU/alu_shift/C86/n27 ), .Z(n17111)
         );
  OAI21_X2 U12354 ( .B1(n17662), .B2(n17306), .A(n16689), .ZN(
        \pipeline/stageE/input1_to_ALU [3]) );
  INV_X2 U12355 ( .A(\pipeline/stageE/input2_to_ALU[0] ), .ZN(n17742) );
  NOR2_X2 U12356 ( .A1(n17387), .A2(n14982), .ZN(n16607) );
  INV_X2 U12357 ( .A(n17741), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[1] ) );
  INV_X4 U12358 ( .A(n17302), .ZN(n17112) );
  INV_X4 U12359 ( .A(n17303), .ZN(n17099) );
  CLKBUF_X1 U12360 ( .A(\pipeline/stageE/EXE_ALU/alu_shift/C48/SH[3] ), .Z(
        n17300) );
  CLKBUF_X1 U12361 ( .A(\pipeline/stageE/EXE_ALU/alu_shift/C48/SH[3] ), .Z(
        n17301) );
  CLKBUF_X1 U12362 ( .A(\pipeline/stageE/EXE_ALU/alu_shift/C48/SH[3] ), .Z(
        n17299) );
  CLKBUF_X1 U12363 ( .A(\pipeline/stageE/EXE_ALU/alu_shift/C48/SH[1] ), .Z(
        n17298) );
  INV_X2 U12364 ( .A(n17739), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[3] ) );
  INV_X2 U12365 ( .A(n13281), .ZN(n17703) );
  AOI21_X1 U12366 ( .B1(n17164), .B2(\pipeline/nextPC_IFID_DEC[25] ), .A(
        n17202), .ZN(\pipeline/stageD/evaluate_jump_target/add_29/n160 ) );
  AOI222_X2 U12367 ( .A1(\pipeline/nextPC_IFID_DEC[1] ), .A2(
        \pipeline/stageD/offset_to_jump_temp [1]), .B1(n17167), .B2(
        \pipeline/nextPC_IFID_DEC[1] ), .C1(
        \pipeline/stageD/evaluate_jump_target/add_29/n214 ), .C2(
        \pipeline/stageD/offset_to_jump_temp [1]), .ZN(n17161) );
  INV_X1 U12368 ( .A(\pipeline/stageE/EXE_ALU/alu_shift/N136 ), .ZN(n17104) );
  INV_X1 U12369 ( .A(\pipeline/stageE/input1_to_ALU [3]), .ZN(n17077) );
  INV_X1 U12370 ( .A(\pipeline/stageE/input1_to_ALU [27]), .ZN(n17078) );
  INV_X1 U12371 ( .A(\pipeline/stageE/input1_to_ALU [17]), .ZN(n17079) );
  INV_X1 U12372 ( .A(\pipeline/stageE/input1_to_ALU [12]), .ZN(n17080) );
  INV_X1 U12373 ( .A(n17074), .ZN(n17081) );
  INV_X1 U12374 ( .A(\pipeline/stageE/input1_to_ALU [11]), .ZN(n17082) );
  INV_X1 U12375 ( .A(\pipeline/stageE/input1_to_ALU [21]), .ZN(n17084) );
  INV_X1 U12376 ( .A(\pipeline/stageE/input1_to_ALU [10]), .ZN(n17085) );
  OAI21_X1 U12377 ( .B1(n17121), .B2(n17320), .A(n16684), .ZN(
        \pipeline/stageE/input1_to_ALU [4]) );
  INV_X1 U12378 ( .A(\pipeline/stageE/input1_to_ALU [26]), .ZN(n17086) );
  INV_X1 U12379 ( .A(\pipeline/stageE/input1_to_ALU [6]), .ZN(n17088) );
  INV_X1 U12380 ( .A(\pipeline/stageE/input1_to_ALU [7]), .ZN(n17089) );
  INV_X1 U12381 ( .A(\pipeline/stageE/input1_to_ALU [9]), .ZN(n17090) );
  INV_X1 U12382 ( .A(n12649), .ZN(n17091) );
  INV_X1 U12383 ( .A(\pipeline/stageE/input1_to_ALU [23]), .ZN(n17092) );
  INV_X1 U12384 ( .A(\pipeline/stageE/input1_to_ALU [28]), .ZN(n17093) );
  INV_X1 U12385 ( .A(\pipeline/stageE/input1_to_ALU [29]), .ZN(n17094) );
  INV_X1 U12386 ( .A(\pipeline/stageE/input1_to_ALU [8]), .ZN(n17095) );
  INV_X1 U12387 ( .A(\pipeline/stageE/input1_to_ALU [18]), .ZN(n17096) );
  NAND2_X2 U12388 ( .A1(n17703), .A2(n17422), .ZN(n17418) );
  BUF_X1 U12389 ( .A(n16591), .Z(n17658) );
  BUF_X1 U12390 ( .A(n16595), .Z(n17654) );
  BUF_X1 U12391 ( .A(n13151), .Z(n17713) );
  INV_X2 U12392 ( .A(n16777), .ZN(n17120) );
  AND2_X1 U12393 ( .A1(n17572), .A2(n17662), .ZN(n16620) );
  BUF_X1 U12394 ( .A(n16592), .Z(n17657) );
  BUF_X1 U12395 ( .A(n16593), .Z(n17656) );
  BUF_X1 U12396 ( .A(n16594), .Z(n17655) );
  BUF_X1 U12397 ( .A(n16596), .Z(n17651) );
  BUF_X1 U12398 ( .A(n16597), .Z(n17650) );
  BUF_X1 U12399 ( .A(n16590), .Z(n17661) );
  NAND2_X2 U12400 ( .A1(n17670), .A2(n13942), .ZN(n17422) );
  BUF_X1 U12401 ( .A(n16617), .Z(n17105) );
  NOR2_X1 U12402 ( .A1(n17012), .A2(n17013), .ZN(n17660) );
  NOR2_X2 U12403 ( .A1(addr_to_dataRam[2]), .A2(n17013), .ZN(n17530) );
  BUF_X2 U12404 ( .A(n13055), .Z(n17098) );
  BUF_X1 U12405 ( .A(n17672), .Z(n17107) );
  NOR2_X1 U12406 ( .A1(\pipeline/stall ), .A2(n15648), .ZN(n17672) );
  INV_X1 U12407 ( .A(n17420), .ZN(n17109) );
  AOI221_X1 U12408 ( .B1(\pipeline/stageE/EXE_ALU/alu_shift/C50/n51 ), .B2(
        \pipeline/stageE/input1_to_ALU [14]), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n167 ), .C2(n17160), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n132 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n43 ) );
  AOI221_X1 U12409 ( .B1(\pipeline/stageE/EXE_ALU/alu_shift/C48/n2 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/A[16] ), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n53 ), .C2(
        \pipeline/stageE/input1_to_ALU [17]), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n151 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n115 ) );
  AOI221_X1 U12410 ( .B1(\pipeline/stageE/EXE_ALU/alu_shift/C50/n51 ), .B2(
        n17160), .C1(\pipeline/stageE/EXE_ALU/alu_shift/C50/n167 ), .C2(
        \pipeline/stageE/input1_to_ALU [12]), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n144 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n63 ) );
  AOI221_X1 U12411 ( .B1(\pipeline/stageE/EXE_ALU/alu_shift/C48/n2 ), .B2(
        \pipeline/stageE/input1_to_ALU [14]), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n53 ), .C2(
        \pipeline/stageE/input1_to_ALU [15]), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n161 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n134 ) );
  AOI221_X1 U12412 ( .B1(n17156), .B2(\pipeline/stageE/input1_to_ALU [6]), 
        .C1(\pipeline/stageE/EXE_ALU/alu_shift/C48/n53 ), .C2(
        \pipeline/stageE/input1_to_ALU [7]), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n170 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n36 ) );
  AOI221_X1 U12413 ( .B1(n17156), .B2(\pipeline/stageE/input1_to_ALU [7]), 
        .C1(\pipeline/stageE/EXE_ALU/alu_shift/C48/n53 ), .C2(
        \pipeline/stageE/input1_to_ALU [8]), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n100 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n32 ) );
  AOI221_X1 U12414 ( .B1(\pipeline/stageE/EXE_ALU/alu_shift/C48/n2 ), .B2(
        \pipeline/stageE/input1_to_ALU [8]), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n53 ), .C2(
        \pipeline/stageE/input1_to_ALU [9]), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n67 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n26 ) );
  AOI221_X1 U12415 ( .B1(n17156), .B2(\pipeline/stageE/input1_to_ALU [9]), 
        .C1(\pipeline/stageE/EXE_ALU/alu_shift/C48/n53 ), .C2(
        \pipeline/stageE/input1_to_ALU [10]), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n54 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n20 ) );
  INV_X2 U12416 ( .A(\pipeline/stall ), .ZN(n15646) );
  NAND2_X1 U12417 ( .A1(n16693), .A2(\pipeline/stageE/input1_to_ALU [1]), .ZN(
        n15049) );
  NAND2_X1 U12418 ( .A1(\pipeline/stageE/EXE_ALU/alu_shift/C48/SH[1] ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n44 ) );
  OAI21_X1 U12419 ( .B1(n17121), .B2(n17362), .A(n16792), .ZN(
        \pipeline/stageE/input1_to_ALU [30]) );
  INV_X1 U12420 ( .A(\pipeline/stageE/input1_to_ALU [14]), .ZN(n17100) );
  INV_X1 U12421 ( .A(\pipeline/stageE/input1_to_ALU [15]), .ZN(n17101) );
  INV_X1 U12422 ( .A(\pipeline/stageE/input1_to_ALU [4]), .ZN(n17102) );
  INV_X1 U12423 ( .A(\pipeline/stageE/input1_to_ALU [1]), .ZN(n17103) );
  NAND2_X1 U12424 ( .A1(n17653), .A2(n17098), .ZN(n16595) );
  BUF_X1 U12425 ( .A(n16617), .Z(n17121) );
  BUF_X1 U12426 ( .A(n17652), .Z(n17653) );
  BUF_X1 U12427 ( .A(n17668), .Z(n17123) );
  NOR2_X1 U12428 ( .A1(n17012), .A2(n17013), .ZN(n16823) );
  BUF_X1 U12429 ( .A(n16817), .Z(n17124) );
  NOR2_X2 U12430 ( .A1(addr_to_dataRam[2]), .A2(n17013), .ZN(n16824) );
  NOR2_X1 U12431 ( .A1(addr_to_dataRam[4]), .A2(n17016), .ZN(n16819) );
  BUF_X1 U12432 ( .A(n16818), .Z(n17125) );
  NOR2_X1 U12433 ( .A1(n17012), .A2(n17013), .ZN(n17659) );
  INV_X1 U12434 ( .A(n16561), .ZN(n17643) );
  BUF_X1 U12435 ( .A(n14964), .Z(n17126) );
  NOR2_X2 U12436 ( .A1(addr_to_dataRam[3]), .A2(n17014), .ZN(n17531) );
  NOR2_X1 U12437 ( .A1(n17155), .A2(read_notWrite), .ZN(n13055) );
  NOR2_X2 U12438 ( .A1(addr_to_dataRam[3]), .A2(n17014), .ZN(n16821) );
  NOR2_X2 U12439 ( .A1(\pipeline/EXE_controls_in_EXEcute [3]), .A2(n15582), 
        .ZN(n17419) );
  BUF_X1 U12440 ( .A(n15903), .Z(n17142) );
  BUF_X1 U12441 ( .A(n15931), .Z(n17145) );
  BUF_X1 U12442 ( .A(n15918), .Z(n17141) );
  BUF_X1 U12443 ( .A(n15905), .Z(n17144) );
  BUF_X1 U12444 ( .A(n15914), .Z(n17136) );
  BUF_X1 U12445 ( .A(n15912), .Z(n17140) );
  BUF_X1 U12446 ( .A(n15930), .Z(n17143) );
  BUF_X1 U12447 ( .A(n15917), .Z(n17139) );
  BUF_X1 U12448 ( .A(n15926), .Z(n17148) );
  BUF_X1 U12449 ( .A(n15927), .Z(n17131) );
  BUF_X1 U12450 ( .A(n15924), .Z(n17128) );
  BUF_X1 U12451 ( .A(n15928), .Z(n17146) );
  BUF_X1 U12452 ( .A(n15925), .Z(n17134) );
  BUF_X1 U12453 ( .A(n15929), .Z(n17147) );
  BUF_X1 U12454 ( .A(n15940), .Z(n17137) );
  BUF_X1 U12455 ( .A(n15935), .Z(n17135) );
  BUF_X1 U12456 ( .A(n15936), .Z(n17132) );
  BUF_X1 U12457 ( .A(n15937), .Z(n17127) );
  BUF_X1 U12458 ( .A(n15906), .Z(n17133) );
  BUF_X1 U12459 ( .A(n15941), .Z(n17138) );
  BUF_X1 U12460 ( .A(n15938), .Z(n17130) );
  BUF_X1 U12461 ( .A(n15939), .Z(n17129) );
  NOR2_X2 U12462 ( .A1(n14860), .A2(n14866), .ZN(n17417) );
  NOR2_X2 U12463 ( .A1(n14864), .A2(n14861), .ZN(n17413) );
  NOR2_X2 U12464 ( .A1(n14865), .A2(n14861), .ZN(n17414) );
  NOR2_X2 U12465 ( .A1(n14863), .A2(n14861), .ZN(n17415) );
  NOR2_X2 U12466 ( .A1(n14860), .A2(n14861), .ZN(n17416) );
  AOI221_X1 U12467 ( .B1(n17304), .B2(
        \pipeline/stageD/offset_jump_sign_ext [22]), .C1(
        \pipeline/stageD/offset_jump_sign_ext [31]), .C2(n17386), .A(n16568), 
        .ZN(n16565) );
  NOR2_X2 U12468 ( .A1(n13281), .A2(\pipeline/WB_controls_in_MEMWB[0] ), .ZN(
        n17370) );
  INV_X1 U12469 ( .A(n13281), .ZN(n17701) );
  INV_X1 U12470 ( .A(n13281), .ZN(n17702) );
  INV_X2 U12471 ( .A(n13281), .ZN(n17704) );
  NOR3_X1 U12472 ( .A1(n17606), .A2(n17605), .A3(n17604), .ZN(n15218) );
  AOI21_X1 U12473 ( .B1(n16646), .B2(n17591), .A(n17592), .ZN(n15368) );
  AND3_X1 U12474 ( .A1(n17588), .A2(n17589), .A3(n17590), .ZN(n15445) );
  BUF_X1 U12475 ( .A(n15600), .Z(n17671) );
  BUF_X1 U12476 ( .A(n15601), .Z(n17673) );
  BUF_X2 U12477 ( .A(n15608), .Z(n17106) );
  BUF_X2 U12478 ( .A(n15610), .Z(n17108) );
  AOI221_X1 U12479 ( .B1(\pipeline/stageE/EXE_ALU/alu_shift/C48/n2 ), .B2(
        \pipeline/stageE/input1_to_ALU [15]), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n53 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/A[16] ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n132 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n99 ) );
  BUF_X1 U12480 ( .A(n15611), .Z(n17674) );
  AOI221_X1 U12481 ( .B1(\pipeline/stageE/EXE_ALU/alu_shift/C48/n2 ), .B2(
        \pipeline/stageE/input1_to_ALU [11]), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n53 ), .C2(
        \pipeline/stageE/input1_to_ALU [12]), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n94 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n4 ) );
  AOI221_X1 U12482 ( .B1(\pipeline/stageE/EXE_ALU/alu_shift/C48/n2 ), .B2(
        \pipeline/stageE/input1_to_ALU [13]), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n53 ), .C2(
        \pipeline/stageE/input1_to_ALU [14]), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n145 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n45 ) );
  AOI221_X1 U12483 ( .B1(\pipeline/stageE/EXE_ALU/alu_shift/C48/n2 ), .B2(
        \pipeline/stageE/input1_to_ALU [12]), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n53 ), .C2(n17160), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n154 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n64 ) );
  AOI221_X1 U12484 ( .B1(\pipeline/stageE/EXE_ALU/alu_shift/C48/n2 ), .B2(
        \pipeline/stageE/input1_to_ALU [10]), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n53 ), .C2(
        \pipeline/stageE/input1_to_ALU [11]), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n157 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n14 ) );
  BUF_X2 U12485 ( .A(\pipeline/stageE/EXE_ALU/alu_shift/C86/n26 ), .Z(n17110)
         );
  NAND2_X2 U12486 ( .A1(\pipeline/stageE/EXE_ALU/alu_shift/C48/SH[1] ), .A2(
        n17742), .ZN(\pipeline/stageE/EXE_ALU/alu_shift/C86/n21 ) );
  NAND2_X2 U12487 ( .A1(\pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[1] ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n23 ) );
  BUF_X2 U12488 ( .A(\pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .Z(n17113) );
  INV_X2 U12489 ( .A(n17081), .ZN(n17114) );
  INV_X1 U12490 ( .A(\pipeline/stageE/input1_to_ALU [25]), .ZN(n17115) );
  INV_X1 U12491 ( .A(\pipeline/stageE/input1_to_ALU [22]), .ZN(n17116) );
  INV_X1 U12492 ( .A(\pipeline/stageE/input1_to_ALU [24]), .ZN(n17117) );
  INV_X1 U12493 ( .A(\pipeline/stageE/input1_to_ALU [20]), .ZN(n17118) );
  INV_X1 U12494 ( .A(\pipeline/stageE/EXE_ALU/alu_shift/N202 ), .ZN(n17119) );
  BUF_X1 U12495 ( .A(n16620), .Z(n17664) );
  BUF_X1 U12496 ( .A(n13103), .Z(n17729) );
  NAND2_X1 U12497 ( .A1(n17530), .A2(n17098), .ZN(n16591) );
  BUF_X1 U12498 ( .A(n16617), .Z(n17662) );
  BUF_X1 U12499 ( .A(n17669), .Z(n17670) );
  BUF_X2 U12500 ( .A(n16619), .Z(n17663) );
  BUF_X2 U12501 ( .A(n16819), .Z(n17122) );
  NOR3_X1 U12502 ( .A1(addr_to_dataRam[4]), .A2(addr_to_dataRam[2]), .A3(
        n17015), .ZN(n17652) );
  NAND2_X2 U12503 ( .A1(\pipeline/stageE/EXE_ALU/add_alu/sCout[0] ), .A2(
        n15573), .ZN(n14968) );
  BUF_X2 U12504 ( .A(n14213), .Z(n17700) );
  BUF_X1 U12505 ( .A(n14246), .Z(n17687) );
  BUF_X2 U12506 ( .A(n14225), .Z(n17698) );
  BUF_X1 U12507 ( .A(n14238), .Z(n17691) );
  BUF_X1 U12508 ( .A(n14250), .Z(n17683) );
  BUF_X1 U12509 ( .A(n14240), .Z(n17689) );
  BUF_X2 U12510 ( .A(n14247), .Z(n17684) );
  BUF_X2 U12511 ( .A(n14239), .Z(n17688) );
  BUF_X1 U12512 ( .A(n14248), .Z(n17685) );
  BUF_X1 U12513 ( .A(n14222), .Z(n17699) );
  BUF_X2 U12514 ( .A(n14244), .Z(n17686) );
  BUF_X1 U12515 ( .A(n14236), .Z(n17693) );
  BUF_X1 U12516 ( .A(n14234), .Z(n17695) );
  BUF_X2 U12517 ( .A(n14227), .Z(n17696) );
  BUF_X2 U12518 ( .A(n14237), .Z(n17690) );
  BUF_X1 U12519 ( .A(n14228), .Z(n17697) );
  BUF_X2 U12520 ( .A(n14233), .Z(n17694) );
  BUF_X2 U12521 ( .A(n14235), .Z(n17692) );
  NOR2_X2 U12522 ( .A1(n16529), .A2(n16531), .ZN(n17392) );
  NOR2_X2 U12523 ( .A1(n16530), .A2(n16534), .ZN(n17390) );
  NOR2_X2 U12524 ( .A1(n16532), .A2(n16534), .ZN(n17389) );
  NOR2_X2 U12525 ( .A1(n16527), .A2(n16534), .ZN(n17388) );
  NOR2_X2 U12526 ( .A1(n16527), .A2(n16528), .ZN(n17391) );
  BUF_X2 U12527 ( .A(n14966), .Z(n17149) );
  BUF_X2 U12528 ( .A(n14965), .Z(n17150) );
  BUF_X2 U12529 ( .A(n14215), .Z(n17151) );
  BUF_X2 U12530 ( .A(n14224), .Z(n17152) );
  BUF_X2 U12531 ( .A(n14245), .Z(n17153) );
  BUF_X2 U12532 ( .A(n14249), .Z(n17154) );
  CLKBUF_X1 U12533 ( .A(\pipeline/Forward_sw1_mux ), .Z(n17744) );
  INV_X1 U12534 ( .A(\pipeline/Forward_sw1_mux ), .ZN(n17743) );
  NOR2_X2 U12535 ( .A1(n16530), .A2(n16534), .ZN(n15913) );
  NOR2_X2 U12536 ( .A1(n16532), .A2(n16534), .ZN(n15915) );
  NOR2_X2 U12537 ( .A1(n16527), .A2(n16528), .ZN(n15901) );
  NOR2_X2 U12538 ( .A1(\pipeline/EXE_controls_in_EXEcute [3]), .A2(n15582), 
        .ZN(n14961) );
  OAI21_X2 U12539 ( .B1(n17105), .B2(n17425), .A(n16793), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N136 ) );
  INV_X1 U12540 ( .A(\pipeline/stageE/EXE_ALU/alu_shift/C48/n46 ), .ZN(n17156)
         );
  NOR2_X2 U12541 ( .A1(n17742), .A2(n17303), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n53 ) );
  NOR2_X2 U12542 ( .A1(n17411), .A2(n15588), .ZN(n14954) );
  INV_X1 U12543 ( .A(n17118), .ZN(n17157) );
  NOR2_X2 U12544 ( .A1(n17074), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[3] ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n1 ) );
  OAI21_X2 U12545 ( .B1(n17662), .B2(n17318), .A(n16678), .ZN(
        \pipeline/stageE/input1_to_ALU [6]) );
  OAI21_X2 U12546 ( .B1(n17121), .B2(n17423), .A(n16637), .ZN(
        \pipeline/stageE/input1_to_ALU [19]) );
  OAI21_X2 U12547 ( .B1(n17105), .B2(n17363), .A(n16734), .ZN(
        \pipeline/stageE/input1_to_ALU [18]) );
  OAI21_X2 U12548 ( .B1(n17105), .B2(n17365), .A(n16770), .ZN(
        \pipeline/stageE/input1_to_ALU [29]) );
  INV_X2 U12549 ( .A(n14981), .ZN(n14952) );
  INV_X1 U12550 ( .A(n17117), .ZN(n17158) );
  OAI21_X2 U12551 ( .B1(n17105), .B2(n17309), .A(n16653), .ZN(
        \pipeline/stageE/input1_to_ALU [14]) );
  OAI21_X2 U12552 ( .B1(n17105), .B2(n17325), .A(n16762), .ZN(
        \pipeline/stageE/input1_to_ALU [27]) );
  OAI21_X2 U12553 ( .B1(n17121), .B2(n17424), .A(n16758), .ZN(
        \pipeline/stageE/input1_to_ALU [26]) );
  OAI21_X2 U12554 ( .B1(n17121), .B2(n17364), .A(n16733), .ZN(
        \pipeline/stageE/input1_to_ALU [15]) );
  OAI21_X2 U12555 ( .B1(n17121), .B2(n17307), .A(n16721), .ZN(
        \pipeline/stageE/input1_to_ALU [10]) );
  OAI21_X2 U12556 ( .B1(n17105), .B2(n17305), .A(n16671), .ZN(
        \pipeline/stageE/input1_to_ALU [9]) );
  INV_X1 U12557 ( .A(n17115), .ZN(n17159) );
  OAI21_X2 U12558 ( .B1(n17105), .B2(n17312), .A(n16766), .ZN(
        \pipeline/stageE/input1_to_ALU [28]) );
  OAI21_X2 U12559 ( .B1(n17121), .B2(n17343), .A(n16713), .ZN(
        \pipeline/stageE/input1_to_ALU [7]) );
  OAI21_X2 U12560 ( .B1(n17121), .B2(n17394), .A(n16720), .ZN(
        \pipeline/stageE/input1_to_ALU [8]) );
  OAI21_X2 U12561 ( .B1(n17121), .B2(n17395), .A(n16660), .ZN(
        \pipeline/stageE/input1_to_ALU [12]) );
  OAI21_X2 U12562 ( .B1(n17105), .B2(n17323), .A(n16645), .ZN(
        \pipeline/stageE/input1_to_ALU [17]) );
  OAI21_X2 U12563 ( .B1(n17105), .B2(n17319), .A(n16725), .ZN(
        \pipeline/stageE/input1_to_ALU [11]) );
  OAI21_X2 U12564 ( .B1(n17121), .B2(n17311), .A(n16749), .ZN(
        \pipeline/stageE/input1_to_ALU [22]) );
  OAI21_X2 U12565 ( .B1(n17121), .B2(n17310), .A(n16742), .ZN(
        \pipeline/stageE/input1_to_ALU [21]) );
  OAI21_X2 U12566 ( .B1(n17105), .B2(n17366), .A(n16753), .ZN(
        \pipeline/stageE/input1_to_ALU [23]) );
  INV_X1 U12567 ( .A(n15425), .ZN(n17160) );
  INV_X4 U12568 ( .A(n17742), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ) );
  NOR4_X2 U12569 ( .A1(\pipeline/stageD/offset_to_jump_temp [10]), .A2(
        \pipeline/stageD/offset_to_jump_temp [9]), .A3(
        \pipeline/stageD/offset_to_jump_temp [7]), .A4(n14174), .ZN(n14005) );
  NOR2_X2 U12570 ( .A1(n16529), .A2(n16531), .ZN(n15907) );
  NOR2_X2 U12571 ( .A1(n16527), .A2(n16534), .ZN(n15916) );
  NOR2_X2 U12572 ( .A1(n17411), .A2(n15588), .ZN(n17677) );
  NOR2_X2 U12573 ( .A1(n17074), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[3] ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n1 ) );
  AND2_X2 U12574 ( .A1(\pipeline/WB_controls_in_MEMWB[0] ), .A2(n17705), .ZN(
        n14135) );
  XNOR2_X1 U12575 ( .A(\pipeline/stageD/evaluate_jump_target/add_29/n138 ), 
        .B(\pipeline/stageD/evaluate_jump_target/add_29/n139 ), .ZN(
        \pipeline/stageD/evaluate_jump_target/N38 ) );
  XNOR2_X1 U12576 ( .A(n17163), .B(
        \pipeline/stageD/evaluate_jump_target/add_29/n201 ), .ZN(
        \pipeline/stageD/evaluate_jump_target/N47 ) );
  XNOR2_X1 U12577 ( .A(\pipeline/stageD/evaluate_jump_target/add_29/n191 ), 
        .B(n17169), .ZN(\pipeline/stageD/evaluate_jump_target/N50 ) );
  XNOR2_X1 U12578 ( .A(\pipeline/stageD/evaluate_jump_target/add_29/n172 ), 
        .B(\pipeline/stageD/evaluate_jump_target/add_29/n175 ), .ZN(
        \pipeline/stageD/evaluate_jump_target/N55 ) );
  XNOR2_X1 U12579 ( .A(\pipeline/stageD/evaluate_jump_target/add_29/n171 ), 
        .B(n17166), .ZN(\pipeline/stageD/evaluate_jump_target/N56 ) );
  XNOR2_X1 U12580 ( .A(\pipeline/stageD/evaluate_jump_target/add_29/n197 ), 
        .B(\pipeline/stageD/evaluate_jump_target/add_29/n196 ), .ZN(
        \pipeline/stageD/evaluate_jump_target/N48 ) );
  XNOR2_X1 U12581 ( .A(\pipeline/stageD/evaluate_jump_target/add_29/n144 ), 
        .B(n17182), .ZN(\pipeline/stageD/evaluate_jump_target/N36 ) );
  XNOR2_X1 U12582 ( .A(\pipeline/stageD/evaluate_jump_target/add_29/n165 ), 
        .B(n17164), .ZN(\pipeline/stageD/evaluate_jump_target/N58 ) );
  XNOR2_X1 U12583 ( .A(n17171), .B(
        \pipeline/stageD/evaluate_jump_target/add_29/n181 ), .ZN(
        \pipeline/stageD/evaluate_jump_target/N53 ) );
  XNOR2_X1 U12584 ( .A(n17162), .B(
        \pipeline/stageD/evaluate_jump_target/add_29/n195 ), .ZN(
        \pipeline/stageD/evaluate_jump_target/N49 ) );
  XNOR2_X1 U12585 ( .A(\pipeline/stageD/evaluate_jump_target/add_29/n177 ), 
        .B(n17179), .ZN(\pipeline/stageD/evaluate_jump_target/N54 ) );
  XNOR2_X1 U12586 ( .A(\pipeline/stageD/evaluate_jump_target/add_29/n126 ), 
        .B(n17175), .ZN(\pipeline/stageD/evaluate_jump_target/N42 ) );
  XNOR2_X1 U12587 ( .A(\pipeline/stageD/evaluate_jump_target/add_29/n132 ), 
        .B(\pipeline/stageD/evaluate_jump_target/add_29/n133 ), .ZN(
        \pipeline/stageD/evaluate_jump_target/N40 ) );
  XNOR2_X1 U12588 ( .A(n17161), .B(
        \pipeline/stageD/evaluate_jump_target/add_29/n150 ), .ZN(
        \pipeline/stageD/evaluate_jump_target/N35 ) );
  XNOR2_X1 U12589 ( .A(n17168), .B(
        \pipeline/stageD/evaluate_jump_target/add_29/n189 ), .ZN(
        \pipeline/stageD/evaluate_jump_target/N51 ) );
  XNOR2_X1 U12590 ( .A(\pipeline/stageD/evaluate_jump_target/add_29/n134 ), 
        .B(\pipeline/stageD/evaluate_jump_target/add_29/n135 ), .ZN(
        \pipeline/stageD/evaluate_jump_target/N39 ) );
  XNOR2_X1 U12591 ( .A(\pipeline/stageD/evaluate_jump_target/add_29/n160 ), 
        .B(\pipeline/stageD/evaluate_jump_target/add_29/n163 ), .ZN(
        \pipeline/stageD/evaluate_jump_target/N59 ) );
  XNOR2_X1 U12592 ( .A(n17173), .B(
        \pipeline/stageD/evaluate_jump_target/add_29/n213 ), .ZN(
        \pipeline/stageD/evaluate_jump_target/N43 ) );
  XNOR2_X1 U12593 ( .A(n17165), .B(
        \pipeline/stageD/evaluate_jump_target/add_29/n169 ), .ZN(
        \pipeline/stageD/evaluate_jump_target/N57 ) );
  NAND2_X1 U12594 ( .A1(net175543), .A2(\pipeline/nextPC_IFID_DEC[0] ), .ZN(
        \pipeline/stageD/evaluate_jump_target/add_29/n183 ) );
  AOI222_X1 U12595 ( .A1(\pipeline/nextPC_IFID_DEC[13] ), .A2(
        \pipeline/stageD/offset_to_jump_temp [13]), .B1(
        \pipeline/nextPC_IFID_DEC[13] ), .B2(
        \pipeline/stageD/evaluate_jump_target/add_29/n202 ), .C1(
        \pipeline/stageD/offset_to_jump_temp [13]), .C2(
        \pipeline/stageD/evaluate_jump_target/add_29/n202 ), .ZN(n17163) );
  XNOR2_X1 U12596 ( .A(n17180), .B(
        \pipeline/stageD/evaluate_jump_target/add_29/n141 ), .ZN(
        \pipeline/stageD/evaluate_jump_target/N37 ) );
  AOI22_X1 U12597 ( .A1(\pipeline/nextPC_IFID_DEC[2] ), .A2(
        \pipeline/stageD/offset_to_jump_temp [2]), .B1(n17404), .B2(n17470), 
        .ZN(\pipeline/stageD/evaluate_jump_target/add_29/n150 ) );
  AOI222_X1 U12598 ( .A1(\pipeline/nextPC_IFID_DEC[23] ), .A2(
        \pipeline/stageD/offset_to_jump_temp [23]), .B1(
        \pipeline/nextPC_IFID_DEC[23] ), .B2(n17166), .C1(
        \pipeline/stageD/offset_to_jump_temp [23]), .C2(n17166), .ZN(n17165)
         );
  AOI222_X1 U12599 ( .A1(\pipeline/nextPC_IFID_DEC[17] ), .A2(
        \pipeline/stageD/offset_to_jump_temp [17]), .B1(
        \pipeline/nextPC_IFID_DEC[17] ), .B2(n17169), .C1(
        \pipeline/stageD/evaluate_jump_target/add_29/n190 ), .C2(
        \pipeline/stageD/offset_to_jump_temp [17]), .ZN(n17168) );
  XNOR2_X1 U12600 ( .A(\pipeline/stageD/evaluate_jump_target/add_29/n185 ), 
        .B(\pipeline/stageD/evaluate_jump_target/add_29/n182 ), .ZN(
        \pipeline/stageD/evaluate_jump_target/N52 ) );
  AOI222_X1 U12601 ( .A1(\pipeline/nextPC_IFID_DEC[19] ), .A2(
        \pipeline/stageD/offset_to_jump_temp [19]), .B1(
        \pipeline/stageD/evaluate_jump_target/add_29/n182 ), .B2(
        \pipeline/nextPC_IFID_DEC[19] ), .C1(
        \pipeline/stageD/evaluate_jump_target/add_29/n182 ), .C2(
        \pipeline/stageD/offset_to_jump_temp [19]), .ZN(n17172) );
  AOI222_X1 U12602 ( .A1(\pipeline/nextPC_IFID_DEC[19] ), .A2(
        \pipeline/stageD/offset_to_jump_temp [19]), .B1(
        \pipeline/nextPC_IFID_DEC[19] ), .B2(
        \pipeline/stageD/evaluate_jump_target/add_29/n182 ), .C1(
        \pipeline/stageD/evaluate_jump_target/add_29/n182 ), .C2(
        \pipeline/stageD/offset_to_jump_temp [19]), .ZN(n17171) );
  AOI222_X1 U12603 ( .A1(\pipeline/stageD/offset_to_jump_temp [9]), .A2(
        \pipeline/nextPC_IFID_DEC[9] ), .B1(
        \pipeline/stageD/offset_to_jump_temp [9]), .B2(n17175), .C1(
        \pipeline/nextPC_IFID_DEC[9] ), .C2(n17175), .ZN(n17173) );
  XNOR2_X1 U12604 ( .A(\pipeline/stageD/evaluate_jump_target/add_29/n128 ), 
        .B(\pipeline/stageD/evaluate_jump_target/add_29/n129 ), .ZN(
        \pipeline/stageD/evaluate_jump_target/N41 ) );
  AOI222_X1 U12605 ( .A1(\pipeline/nextPC_IFID_DEC[11] ), .A2(
        \pipeline/stageD/offset_to_jump_temp [11]), .B1(
        \pipeline/stageD/evaluate_jump_target/add_29/n208 ), .B2(
        \pipeline/nextPC_IFID_DEC[11] ), .C1(
        \pipeline/stageD/evaluate_jump_target/add_29/n208 ), .C2(
        \pipeline/stageD/offset_to_jump_temp [11]), .ZN(n17178) );
  XNOR2_X1 U12606 ( .A(\pipeline/stageD/evaluate_jump_target/add_29/n203 ), 
        .B(\pipeline/stageD/evaluate_jump_target/add_29/n202 ), .ZN(
        \pipeline/stageD/evaluate_jump_target/N46 ) );
  AOI222_X1 U12607 ( .A1(\pipeline/nextPC_IFID_DEC[3] ), .A2(
        \pipeline/stageD/offset_to_jump_temp [3]), .B1(
        \pipeline/nextPC_IFID_DEC[3] ), .B2(n17182), .C1(
        \pipeline/stageD/offset_to_jump_temp [3]), .C2(n17182), .ZN(n17180) );
  AOI222_X1 U12608 ( .A1(n17161), .A2(n17470), .B1(
        \pipeline/stageD/evaluate_jump_target/add_29/n149 ), .B2(n17404), .C1(
        n17470), .C2(n17404), .ZN(
        \pipeline/stageD/evaluate_jump_target/add_29/n145 ) );
  NAND3_X1 U12609 ( .A1(n17186), .A2(n17185), .A3(n17184), .ZN(n17188) );
  XNOR2_X1 U12610 ( .A(n17192), .B(n17191), .ZN(
        \pipeline/stageD/evaluate_jump_target/N62 ) );
  NAND2_X1 U12611 ( .A1(n17190), .A2(n17189), .ZN(n17192) );
  AOI21_X1 U12612 ( .B1(n17201), .B2(n17451), .A(n17200), .ZN(n17202) );
  NAND2_X1 U12613 ( .A1(n17166), .A2(\pipeline/stageD/offset_to_jump_temp [23]), .ZN(n17195) );
  NAND2_X1 U12614 ( .A1(\pipeline/stageD/evaluate_jump_target/add_29/n170 ), 
        .A2(\pipeline/stageD/offset_to_jump_temp [23]), .ZN(n17194) );
  NAND3_X1 U12615 ( .A1(n17196), .A2(
        \pipeline/stageD/evaluate_jump_target/add_29/n168 ), .A3(n17194), .ZN(
        n17199) );
  NAND3_X1 U12616 ( .A1(n17196), .A2(n17465), .A3(n17195), .ZN(n17198) );
  NAND3_X1 U12617 ( .A1(n17198), .A2(n17199), .A3(n17197), .ZN(n17201) );
  NAND2_X1 U12618 ( .A1(n17208), .A2(n17465), .ZN(n17207) );
  NAND2_X1 U12619 ( .A1(\pipeline/stageD/evaluate_jump_target/add_29/n168 ), 
        .A2(n17208), .ZN(n17209) );
  OAI21_X1 U12620 ( .B1(n17464), .B2(
        \pipeline/stageD/evaluate_jump_target/add_29/n174 ), .A(
        \pipeline/stageD/evaluate_jump_target/add_29/n172 ), .ZN(n17214) );
  AOI21_X1 U12621 ( .B1(n17219), .B2(n17448), .A(n17218), .ZN(n17220) );
  NAND2_X1 U12622 ( .A1(\pipeline/stageD/evaluate_jump_target/add_29/n178 ), 
        .A2(\pipeline/stageD/evaluate_jump_target/add_29/n180 ), .ZN(n17217)
         );
  NAND2_X1 U12623 ( .A1(n17172), .A2(n17463), .ZN(n17216) );
  NAND3_X1 U12624 ( .A1(n17216), .A2(n17217), .A3(n17215), .ZN(n17219) );
  AOI222_X1 U12625 ( .A1(\pipeline/nextPC_IFID_DEC[19] ), .A2(
        \pipeline/stageD/offset_to_jump_temp [19]), .B1(
        \pipeline/stageD/evaluate_jump_target/add_29/n182 ), .B2(
        \pipeline/nextPC_IFID_DEC[19] ), .C1(
        \pipeline/stageD/evaluate_jump_target/add_29/n182 ), .C2(
        \pipeline/stageD/offset_to_jump_temp [19]), .ZN(
        \pipeline/stageD/evaluate_jump_target/add_29/n178 ) );
  NAND2_X1 U12626 ( .A1(\pipeline/stageD/evaluate_jump_target/add_29/n190 ), 
        .A2(\pipeline/stageD/offset_to_jump_temp [17]), .ZN(n17222) );
  OAI211_X1 U12627 ( .C1(n17294), .C2(n17290), .A(n17223), .B(n17222), .ZN(
        n17225) );
  NAND2_X1 U12628 ( .A1(\pipeline/stageD/evaluate_jump_target/add_29/n190 ), 
        .A2(\pipeline/nextPC_IFID_DEC[17] ), .ZN(n17223) );
  OAI21_X1 U12629 ( .B1(\pipeline/stageD/evaluate_jump_target/add_29/n174 ), 
        .B2(n17464), .A(\pipeline/stageD/evaluate_jump_target/add_29/n172 ), 
        .ZN(n17227) );
  NAND2_X1 U12630 ( .A1(\pipeline/stageD/evaluate_jump_target/add_29/n196 ), 
        .A2(\pipeline/stageD/offset_to_jump_temp [15]), .ZN(n17230) );
  OAI21_X1 U12631 ( .B1(\pipeline/stageD/evaluate_jump_target/add_29/n196 ), 
        .B2(\pipeline/stageD/offset_to_jump_temp [15]), .A(
        \pipeline/nextPC_IFID_DEC[15] ), .ZN(n17231) );
  NAND2_X1 U12632 ( .A1(\pipeline/stageD/evaluate_jump_target/add_29/n196 ), 
        .A2(\pipeline/stageD/offset_to_jump_temp [15]), .ZN(n17232) );
  OAI21_X1 U12633 ( .B1(\pipeline/stageD/evaluate_jump_target/add_29/n196 ), 
        .B2(\pipeline/stageD/offset_to_jump_temp [15]), .A(
        \pipeline/nextPC_IFID_DEC[15] ), .ZN(n17233) );
  NAND2_X1 U12634 ( .A1(\pipeline/stageD/evaluate_jump_target/add_29/n178 ), 
        .A2(\pipeline/stageD/evaluate_jump_target/add_29/n180 ), .ZN(n17236)
         );
  NAND2_X1 U12635 ( .A1(n17172), .A2(n17463), .ZN(n17235) );
  NAND2_X1 U12636 ( .A1(\pipeline/stageD/evaluate_jump_target/add_29/n202 ), 
        .A2(\pipeline/stageD/offset_to_jump_temp [13]), .ZN(n17238) );
  OAI211_X1 U12637 ( .C1(n17292), .C2(n17288), .A(n17238), .B(n17239), .ZN(
        n17241) );
  NAND2_X1 U12638 ( .A1(\pipeline/stageD/evaluate_jump_target/add_29/n202 ), 
        .A2(\pipeline/nextPC_IFID_DEC[13] ), .ZN(n17239) );
  NAND2_X1 U12639 ( .A1(\pipeline/stageD/evaluate_jump_target/add_29/n208 ), 
        .A2(\pipeline/stageD/offset_to_jump_temp [11]), .ZN(n17243) );
  OAI211_X1 U12640 ( .C1(n17293), .C2(n17289), .A(n17243), .B(n17244), .ZN(
        n17246) );
  NAND2_X1 U12641 ( .A1(\pipeline/stageD/evaluate_jump_target/add_29/n208 ), 
        .A2(\pipeline/nextPC_IFID_DEC[11] ), .ZN(n17244) );
  OAI21_X1 U12642 ( .B1(n17457), .B2(n17428), .A(
        \pipeline/stageD/evaluate_jump_target/add_29/n128 ), .ZN(n17251) );
  OAI22_X1 U12643 ( .A1(n17255), .A2(n17254), .B1(
        \pipeline/nextPC_IFID_DEC[10] ), .B2(
        \pipeline/stageD/offset_to_jump_temp [10]), .ZN(n17256) );
  NAND2_X1 U12644 ( .A1(n17176), .A2(\pipeline/nextPC_IFID_DEC[9] ), .ZN(
        n17248) );
  AOI21_X1 U12645 ( .B1(n17176), .B2(\pipeline/stageD/offset_to_jump_temp [9]), 
        .A(n17247), .ZN(n17249) );
  NAND3_X1 U12646 ( .A1(n17251), .A2(\pipeline/nextPC_IFID_DEC[9] ), .A3(
        n17250), .ZN(n17253) );
  NAND3_X1 U12647 ( .A1(n17253), .A2(n17440), .A3(n17252), .ZN(n17254) );
  OAI21_X1 U12648 ( .B1(n17428), .B2(n17457), .A(
        \pipeline/stageD/evaluate_jump_target/add_29/n128 ), .ZN(n17259) );
  NAND2_X1 U12649 ( .A1(\pipeline/stageD/evaluate_jump_target/add_29/n133 ), 
        .A2(\pipeline/stageD/offset_to_jump_temp [7]), .ZN(n17260) );
  OAI21_X1 U12650 ( .B1(\pipeline/stageD/evaluate_jump_target/add_29/n133 ), 
        .B2(\pipeline/stageD/offset_to_jump_temp [7]), .A(
        \pipeline/nextPC_IFID_DEC[7] ), .ZN(n17261) );
  OAI21_X1 U12651 ( .B1(n17361), .B2(n17456), .A(
        \pipeline/stageD/evaluate_jump_target/add_29/n134 ), .ZN(n17263) );
  NAND2_X1 U12652 ( .A1(\pipeline/nextPC_IFID_DEC[5] ), .A2(
        \pipeline/stageD/offset_to_jump_temp [5]), .ZN(n17266) );
  NAND2_X1 U12653 ( .A1(\pipeline/nextPC_IFID_DEC[5] ), .A2(
        \pipeline/stageD/evaluate_jump_target/add_29/n139 ), .ZN(n17265) );
  NAND2_X1 U12654 ( .A1(\pipeline/stageD/evaluate_jump_target/add_29/n139 ), 
        .A2(\pipeline/stageD/offset_to_jump_temp [5]), .ZN(n17264) );
  NAND2_X1 U12655 ( .A1(\pipeline/stageD/evaluate_jump_target/add_29/n145 ), 
        .A2(\pipeline/stageD/offset_to_jump_temp [3]), .ZN(n17269) );
  AOI21_X1 U12656 ( .B1(\pipeline/stageD/evaluate_jump_target/add_29/n145 ), 
        .B2(\pipeline/nextPC_IFID_DEC[3] ), .A(n17291), .ZN(n17270) );
  NAND2_X1 U12657 ( .A1(n17181), .A2(\pipeline/stageD/offset_to_jump_temp [3]), 
        .ZN(n17267) );
  AOI21_X1 U12658 ( .B1(n17181), .B2(\pipeline/nextPC_IFID_DEC[3] ), .A(n17291), .ZN(n17268) );
  NAND3_X1 U12659 ( .A1(n17268), .A2(n17455), .A3(n17267), .ZN(n17273) );
  NAND3_X1 U12660 ( .A1(n17270), .A2(n17412), .A3(n17269), .ZN(n17271) );
  AOI222_X1 U12661 ( .A1(\pipeline/nextPC_IFID_DEC[1] ), .A2(
        \pipeline/stageD/offset_to_jump_temp [1]), .B1(n17167), .B2(
        \pipeline/nextPC_IFID_DEC[1] ), .C1(
        \pipeline/stageD/evaluate_jump_target/add_29/n214 ), .C2(
        \pipeline/stageD/offset_to_jump_temp [1]), .ZN(n17274) );
  NAND2_X1 U12662 ( .A1(net175543), .A2(\pipeline/nextPC_IFID_DEC[0] ), .ZN(
        n17275) );
  AOI21_X1 U12663 ( .B1(n17406), .B2(n17275), .A(n17446), .ZN(n17277) );
  XNOR2_X1 U12664 ( .A(n17188), .B(n17187), .ZN(
        \pipeline/stageD/evaluate_jump_target/N63 ) );
  NAND3_X1 U12665 ( .A1(n17278), .A2(n17279), .A3(n17287), .ZN(n17185) );
  NAND2_X1 U12666 ( .A1(n17281), .A2(n17200), .ZN(n17278) );
  NAND2_X1 U12667 ( .A1(n17280), .A2(n17286), .ZN(n17190) );
  XNOR2_X1 U12668 ( .A(n17280), .B(
        \pipeline/stageD/evaluate_jump_target/add_29/n157 ), .ZN(
        \pipeline/stageD/evaluate_jump_target/N61 ) );
  NAND2_X1 U12669 ( .A1(n17281), .A2(n17467), .ZN(n17279) );
  NAND2_X1 U12670 ( .A1(n17283), .A2(\pipeline/stageD/offset_to_jump_temp [30]), .ZN(n17193) );
  XNOR2_X1 U12671 ( .A(n17283), .B(
        \pipeline/stageD/evaluate_jump_target/add_29/n159 ), .ZN(
        \pipeline/stageD/evaluate_jump_target/N60 ) );
  OAI21_X1 U12672 ( .B1(n17283), .B2(\pipeline/stageD/offset_to_jump_temp [30]), .A(\pipeline/nextPC_IFID_DEC[27] ), .ZN(n17282) );
  NAND2_X1 U12673 ( .A1(\pipeline/stageD/offset_to_jump_temp [17]), .A2(
        \pipeline/nextPC_IFID_DEC[17] ), .ZN(n17221) );
  NAND2_X1 U12674 ( .A1(\pipeline/stageD/offset_to_jump_temp [13]), .A2(
        \pipeline/nextPC_IFID_DEC[13] ), .ZN(n17237) );
  NAND2_X1 U12675 ( .A1(\pipeline/stageD/offset_to_jump_temp [11]), .A2(
        \pipeline/nextPC_IFID_DEC[11] ), .ZN(n17242) );
  NAND2_X1 U12676 ( .A1(n17412), .A2(n17455), .ZN(n17272) );
  NAND2_X1 U12677 ( .A1(n17361), .A2(n17456), .ZN(n17262) );
  NAND2_X1 U12678 ( .A1(n17428), .A2(n17457), .ZN(n17258) );
  NAND2_X1 U12679 ( .A1(\pipeline/stageD/offset_to_jump_temp [9]), .A2(
        \pipeline/nextPC_IFID_DEC[9] ), .ZN(n17252) );
  NAND2_X1 U12680 ( .A1(n17458), .A2(n17252), .ZN(n17247) );
  NAND2_X1 U12681 ( .A1(n17428), .A2(n17457), .ZN(n17250) );
  NAND2_X1 U12682 ( .A1(n17444), .A2(n17459), .ZN(n17245) );
  NAND2_X1 U12683 ( .A1(n17445), .A2(n17460), .ZN(n17240) );
  NAND2_X1 U12684 ( .A1(\pipeline/stageD/evaluate_jump_target/add_29/n188 ), 
        .A2(n17462), .ZN(n17224) );
  NAND2_X1 U12685 ( .A1(\pipeline/stageD/evaluate_jump_target/add_29/n180 ), 
        .A2(n17463), .ZN(n17234) );
  NAND2_X1 U12686 ( .A1(\pipeline/stageD/evaluate_jump_target/add_29/n180 ), 
        .A2(n17463), .ZN(n17215) );
  NAND2_X1 U12687 ( .A1(\pipeline/stageD/evaluate_jump_target/add_29/n174 ), 
        .A2(n17464), .ZN(n17213) );
  NAND2_X1 U12688 ( .A1(\pipeline/stageD/offset_to_jump_temp [23]), .A2(
        \pipeline/nextPC_IFID_DEC[23] ), .ZN(n17208) );
  NAND2_X1 U12689 ( .A1(\pipeline/stageD/evaluate_jump_target/add_29/n174 ), 
        .A2(n17464), .ZN(n17226) );
  NAND2_X1 U12690 ( .A1(\pipeline/stageD/evaluate_jump_target/add_29/n168 ), 
        .A2(n17465), .ZN(n17210) );
  NAND2_X1 U12691 ( .A1(\pipeline/stageD/evaluate_jump_target/add_29/n168 ), 
        .A2(n17465), .ZN(n17197) );
  NAND2_X1 U12692 ( .A1(n17200), .A2(n17467), .ZN(n17183) );
  NAND2_X1 U12693 ( .A1(\pipeline/stageD/offset_to_jump_temp [30]), .A2(
        \pipeline/nextPC_IFID_DEC[29] ), .ZN(n17184) );
  XNOR2_X1 U12694 ( .A(\pipeline/stageD/offset_to_jump_temp [30]), .B(
        \pipeline/nextPC_IFID_DEC[30] ), .ZN(n17187) );
  NAND2_X1 U12695 ( .A1(n17200), .A2(n17467), .ZN(n17189) );
  XNOR2_X1 U12696 ( .A(\pipeline/stageD/offset_to_jump_temp [30]), .B(n17452), 
        .ZN(n17191) );
  INV_X1 U12697 ( .A(\pipeline/stageD/evaluate_jump_target/add_29/n190 ), .ZN(
        n17170) );
  AND2_X1 U12698 ( .A1(\pipeline/stageD/evaluate_jump_target/add_29/n188 ), 
        .A2(n17221), .ZN(n17294) );
  AND2_X1 U12699 ( .A1(n17221), .A2(n17462), .ZN(n17290) );
  AND2_X1 U12700 ( .A1(n17445), .A2(n17237), .ZN(n17292) );
  AND2_X1 U12701 ( .A1(n17460), .A2(n17237), .ZN(n17288) );
  AND2_X1 U12702 ( .A1(n17444), .A2(n17242), .ZN(n17293) );
  AND2_X1 U12703 ( .A1(n17459), .A2(n17242), .ZN(n17289) );
  AND2_X1 U12704 ( .A1(net175543), .A2(\pipeline/nextPC_IFID_DEC[0] ), .ZN(
        n17167) );
  AND2_X1 U12705 ( .A1(net175543), .A2(\pipeline/nextPC_IFID_DEC[0] ), .ZN(
        \pipeline/stageD/evaluate_jump_target/add_29/n214 ) );
  NOR2_X1 U12706 ( .A1(n17406), .A2(n17275), .ZN(n17276) );
  NOR2_X1 U12707 ( .A1(n17277), .A2(n17276), .ZN(
        \pipeline/stageD/evaluate_jump_target/add_29/n149 ) );
  AND2_X1 U12708 ( .A1(\pipeline/stageD/offset_to_jump_temp [3]), .A2(
        \pipeline/nextPC_IFID_DEC[3] ), .ZN(n17291) );
  AND3_X1 U12709 ( .A1(n17266), .A2(n17265), .A3(n17264), .ZN(
        \pipeline/stageD/evaluate_jump_target/add_29/n134 ) );
  AND2_X1 U12710 ( .A1(n17259), .A2(n17258), .ZN(n17176) );
  AND2_X1 U12711 ( .A1(n17249), .A2(n17248), .ZN(n17257) );
  AND2_X1 U12712 ( .A1(n17177), .A2(\pipeline/stageD/offset_to_jump_temp [9]), 
        .ZN(n17255) );
  AND3_X1 U12713 ( .A1(n17231), .A2(
        \pipeline/stageD/evaluate_jump_target/add_29/n194 ), .A3(n17230), .ZN(
        n17229) );
  AND2_X1 U12714 ( .A1(\pipeline/stageD/evaluate_jump_target/add_29/n194 ), 
        .A2(n17461), .ZN(n17228) );
  AND3_X1 U12715 ( .A1(n17236), .A2(n17235), .A3(n17234), .ZN(n17179) );
  INV_X1 U12716 ( .A(\pipeline/stageD/offset_to_jump_temp [21]), .ZN(n17218)
         );
  AND2_X1 U12717 ( .A1(n17166), .A2(\pipeline/stageD/offset_to_jump_temp [23]), 
        .ZN(n17203) );
  AND2_X1 U12718 ( .A1(n17166), .A2(\pipeline/nextPC_IFID_DEC[23] ), .ZN(
        n17204) );
  OR3_X1 U12719 ( .A1(n17203), .A2(n17204), .A3(n17207), .ZN(n17212) );
  AND2_X1 U12720 ( .A1(n17227), .A2(n17226), .ZN(
        \pipeline/stageD/evaluate_jump_target/add_29/n170 ) );
  AND2_X1 U12721 ( .A1(\pipeline/stageD/evaluate_jump_target/add_29/n170 ), 
        .A2(\pipeline/nextPC_IFID_DEC[23] ), .ZN(n17205) );
  AND2_X1 U12722 ( .A1(\pipeline/stageD/evaluate_jump_target/add_29/n170 ), 
        .A2(\pipeline/stageD/offset_to_jump_temp [23]), .ZN(n17206) );
  OR3_X1 U12723 ( .A1(n17205), .A2(n17206), .A3(n17209), .ZN(n17211) );
  AND3_X1 U12724 ( .A1(n17212), .A2(n17211), .A3(n17210), .ZN(n17164) );
  INV_X1 U12725 ( .A(\pipeline/stageD/offset_to_jump_temp [30]), .ZN(n17200)
         );
  OR2_X1 U12726 ( .A1(n17200), .A2(n17466), .ZN(n17285) );
  AND2_X1 U12727 ( .A1(n17200), .A2(n17466), .ZN(n17284) );
  AND2_X1 U12728 ( .A1(n17282), .A2(n17193), .ZN(n17281) );
  AND2_X1 U12729 ( .A1(n17183), .A2(\pipeline/stageD/offset_to_jump_temp [30]), 
        .ZN(n17287) );
  AND2_X1 U12730 ( .A1(n17282), .A2(n17193), .ZN(n17280) );
  OR2_X1 U12731 ( .A1(n17200), .A2(n17467), .ZN(n17286) );
  INV_X1 U12732 ( .A(n17170), .ZN(n17169) );
  CLKBUF_X1 U12733 ( .A(\pipeline/stageD/evaluate_jump_target/add_29/n208 ), 
        .Z(n17174) );
  CLKBUF_X1 U12734 ( .A(n17177), .Z(n17175) );
  CLKBUF_X1 U12735 ( .A(n17181), .Z(n17182) );
  AOI222_X2 U12736 ( .A1(n17274), .A2(n17470), .B1(
        \pipeline/stageD/evaluate_jump_target/add_29/n149 ), .B2(n17404), .C1(
        n17470), .C2(n17404), .ZN(n17181) );
  NOR2_X2 U12737 ( .A1(n17257), .A2(n17256), .ZN(
        \pipeline/stageD/evaluate_jump_target/add_29/n208 ) );
  AND2_X2 U12738 ( .A1(n17225), .A2(n17224), .ZN(
        \pipeline/stageD/evaluate_jump_target/add_29/n182 ) );
  AND2_X2 U12739 ( .A1(n17214), .A2(n17213), .ZN(n17166) );
  AND2_X2 U12740 ( .A1(n17241), .A2(n17240), .ZN(
        \pipeline/stageD/evaluate_jump_target/add_29/n196 ) );
  AOI21_X1 U12741 ( .B1(\pipeline/stageD/evaluate_jump_target/add_29/n160 ), 
        .B2(n17285), .A(n17284), .ZN(n17283) );
  AND2_X2 U12742 ( .A1(n17246), .A2(n17245), .ZN(
        \pipeline/stageD/evaluate_jump_target/add_29/n202 ) );
  AND3_X2 U12743 ( .A1(n17273), .A2(n17272), .A3(n17271), .ZN(
        \pipeline/stageD/evaluate_jump_target/add_29/n139 ) );
  AOI21_X2 U12744 ( .B1(n17179), .B2(\pipeline/nextPC_IFID_DEC[21] ), .A(
        n17220), .ZN(\pipeline/stageD/evaluate_jump_target/add_29/n172 ) );
  AOI211_X2 U12745 ( .C1(n17162), .C2(n17461), .A(n17229), .B(n17228), .ZN(
        \pipeline/stageD/evaluate_jump_target/add_29/n190 ) );
  AND2_X2 U12746 ( .A1(n17261), .A2(n17260), .ZN(
        \pipeline/stageD/evaluate_jump_target/add_29/n128 ) );
  OR2_X1 U12747 ( .A1(n17428), .A2(n17457), .ZN(n17295) );
  AND2_X1 U12748 ( .A1(\pipeline/stageE/EXE_ALU/alu_shift/N202 ), .A2(n17742), 
        .ZN(\pipeline/stageE/EXE_ALU/alu_shift/C88/ML_int[1][0] ) );
  NAND2_X1 U12749 ( .A1(\pipeline/stageE/EXE_ALU/alu_shift/C48/SH[1] ), .A2(
        n17742), .ZN(\pipeline/stageE/EXE_ALU/alu_shift/C50/n46 ) );
  NOR2_X1 U12750 ( .A1(\pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[1] ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n50 ) );
  NOR2_X1 U12751 ( .A1(n17742), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[1] ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n49 ) );
  NOR2_X1 U12752 ( .A1(n17739), .A2(n17074), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n76 ) );
  AOI22_X1 U12753 ( .A1(\pipeline/stageE/input1_to_ALU [1]), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n26 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/N202 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n27 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n151 ) );
  NOR2_X1 U12754 ( .A1(n17081), .A2(n17296), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n73 ) );
  INV_X1 U12755 ( .A(\pipeline/stageE/EXE_ALU/alu_shift/C50/n46 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n167 ) );
  INV_X1 U12756 ( .A(n17739), .ZN(n17296) );
  INV_X1 U12757 ( .A(n17112), .ZN(n17297) );
  INV_X1 U12758 ( .A(\pipeline/stageE/EXE_ALU/alu_shift/C50/n124 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n72 ) );
  AND2_X1 U12759 ( .A1(n17074), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n148 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C50/n10 ) );
  AND2_X1 U12760 ( .A1(\pipeline/stageE/EXE_ALU/alu_shift/C50/n148 ), .A2(
        n17081), .ZN(\pipeline/stageE/EXE_ALU/alu_shift/C50/n8 ) );
  NOR2_X1 U12761 ( .A1(\pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[1] ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n27 ) );
  NOR2_X1 U12762 ( .A1(n17742), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[1] ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n26 ) );
  AOI222_X1 U12763 ( .A1(n17111), .A2(n12649), .B1(
        \pipeline/stageE/input1_to_ALU [1]), .B2(n17110), .C1(
        \pipeline/stageE/EXE_ALU/alu_shift/N202 ), .C2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[1] ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n170 ) );
  NAND2_X1 U12764 ( .A1(\pipeline/stageE/EXE_ALU/alu_shift/C48/SH[3] ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/N202 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n104 ) );
  NAND2_X1 U12765 ( .A1(\pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/N202 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n4 ) );
  INV_X1 U12766 ( .A(\pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ), .ZN(
        n17302) );
  AND2_X1 U12767 ( .A1(n17074), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[3] ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C86/n136 ) );
  AND2_X1 U12768 ( .A1(\pipeline/stageE/EXE_ALU/alu_shift/C86/n131 ), .A2(
        n17074), .ZN(\pipeline/stageE/EXE_ALU/alu_shift/C86/n15 ) );
  AND2_X1 U12769 ( .A1(\pipeline/stageE/EXE_ALU/alu_shift/C86/n131 ), .A2(
        n17081), .ZN(\pipeline/stageE/EXE_ALU/alu_shift/C86/n19 ) );
  AOI22_X1 U12770 ( .A1(\pipeline/stageE/input1_to_ALU [1]), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n51 ), .B1(
        \pipeline/stageE/EXE_ALU/alu_shift/N202 ), .B2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n52 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n160 ) );
  INV_X1 U12771 ( .A(\pipeline/stageE/EXE_ALU/alu_shift/C48/SH[1] ), .ZN(
        n17303) );
  NOR2_X1 U12772 ( .A1(n17303), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n2 ) );
  AND2_X1 U12773 ( .A1(n17074), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[3] ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n105 ) );
  AND2_X1 U12774 ( .A1(n17074), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n158 ), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/n12 ) );
  AND2_X1 U12775 ( .A1(\pipeline/stageE/EXE_ALU/alu_shift/C48/n158 ), .A2(
        n17081), .ZN(\pipeline/stageE/EXE_ALU/alu_shift/C48/n10 ) );
  OAI21_X1 U12776 ( .B1(n15218), .B2(n15220), .A(n15221), .ZN(n15205) );
  INV_X4 U12777 ( .A(n17737), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[4] ) );
  CLKBUF_X1 U12778 ( .A(n13172), .Z(n17706) );
  CLKBUF_X1 U12779 ( .A(n13166), .Z(n17708) );
  CLKBUF_X1 U12780 ( .A(n13160), .Z(n17710) );
  CLKBUF_X1 U12781 ( .A(n13154), .Z(n17712) );
  CLKBUF_X1 U12782 ( .A(n13148), .Z(n17714) );
  CLKBUF_X1 U12783 ( .A(n13142), .Z(n17716) );
  CLKBUF_X1 U12784 ( .A(n13136), .Z(n17718) );
  CLKBUF_X1 U12785 ( .A(n13130), .Z(n17720) );
  CLKBUF_X1 U12786 ( .A(n13124), .Z(n17722) );
  CLKBUF_X1 U12787 ( .A(n13118), .Z(n17724) );
  CLKBUF_X1 U12788 ( .A(n13112), .Z(n17726) );
  CLKBUF_X1 U12789 ( .A(n13106), .Z(n17728) );
  CLKBUF_X1 U12790 ( .A(n13169), .Z(n17707) );
  CLKBUF_X1 U12791 ( .A(n13163), .Z(n17709) );
  CLKBUF_X1 U12792 ( .A(n13157), .Z(n17711) );
  CLKBUF_X1 U12793 ( .A(n13145), .Z(n17715) );
  CLKBUF_X1 U12794 ( .A(n13139), .Z(n17717) );
  CLKBUF_X1 U12795 ( .A(n13133), .Z(n17719) );
  CLKBUF_X1 U12796 ( .A(n13127), .Z(n17721) );
  CLKBUF_X1 U12797 ( .A(n13121), .Z(n17723) );
  CLKBUF_X1 U12798 ( .A(n13115), .Z(n17725) );
  CLKBUF_X1 U12799 ( .A(n13109), .Z(n17727) );
  CLKBUF_X1 U12800 ( .A(n13097), .Z(n17731) );
  CLKBUF_X1 U12801 ( .A(n13082), .Z(n17736) );
  CLKBUF_X1 U12802 ( .A(n13088), .Z(n17734) );
  CLKBUF_X1 U12803 ( .A(n13094), .Z(n17732) );
  CLKBUF_X1 U12804 ( .A(n13085), .Z(n17735) );
  CLKBUF_X1 U12805 ( .A(n13100), .Z(n17730) );
  CLKBUF_X1 U12806 ( .A(n13091), .Z(n17733) );
  INV_X1 U12807 ( .A(n15116), .ZN(n13184) );
  INV_X1 U12808 ( .A(n15120), .ZN(n13178) );
  INV_X1 U12809 ( .A(n15104), .ZN(n13202) );
  INV_X1 U12810 ( .A(n15112), .ZN(n13190) );
  INV_X1 U12811 ( .A(n15114), .ZN(n13187) );
  INV_X1 U12812 ( .A(n15102), .ZN(n13205) );
  INV_X1 U12813 ( .A(n15108), .ZN(n13196) );
  INV_X1 U12814 ( .A(n15110), .ZN(n13193) );
  INV_X1 U12815 ( .A(n15118), .ZN(n13181) );
  INV_X1 U12816 ( .A(n15084), .ZN(n13232) );
  INV_X1 U12817 ( .A(n15122), .ZN(n13175) );
  INV_X1 U12818 ( .A(n15096), .ZN(n13214) );
  INV_X1 U12819 ( .A(n15092), .ZN(n13220) );
  INV_X1 U12820 ( .A(n15088), .ZN(n13226) );
  INV_X1 U12821 ( .A(n15106), .ZN(n13199) );
  INV_X1 U12822 ( .A(n15064), .ZN(n13262) );
  INV_X1 U12823 ( .A(n15080), .ZN(n13238) );
  INV_X1 U12824 ( .A(n15094), .ZN(n13217) );
  INV_X1 U12825 ( .A(n15076), .ZN(n13244) );
  INV_X1 U12826 ( .A(n15090), .ZN(n13223) );
  INV_X1 U12827 ( .A(n15072), .ZN(n13250) );
  INV_X1 U12828 ( .A(n15082), .ZN(n13235) );
  INV_X1 U12829 ( .A(n15068), .ZN(n13256) );
  INV_X1 U12830 ( .A(n14988), .ZN(n13268) );
  INV_X1 U12831 ( .A(n15062), .ZN(n13265) );
  INV_X1 U12832 ( .A(n15100), .ZN(n13208) );
  INV_X1 U12833 ( .A(n15086), .ZN(n13229) );
  INV_X1 U12834 ( .A(n15074), .ZN(n13247) );
  INV_X1 U12835 ( .A(n15098), .ZN(n13211) );
  INV_X1 U12836 ( .A(n15078), .ZN(n13241) );
  INV_X1 U12837 ( .A(n15066), .ZN(n13259) );
  INV_X1 U12838 ( .A(n15070), .ZN(n13253) );
  INV_X1 U12839 ( .A(n17420), .ZN(n17682) );
  AND2_X1 U12840 ( .A1(n14167), .A2(n14947), .ZN(n17420) );
  AND2_X1 U12841 ( .A1(\pipeline/EXE_controls_in_IDEX[8] ), .A2(
        \pipeline/IDEX_Stage/N181 ), .ZN(\pipeline/IDEX_Stage/N197 ) );
  INV_X1 U12842 ( .A(n15621), .ZN(n3987) );
  AND3_X1 U12843 ( .A1(n17625), .A2(n17626), .A3(n17627), .ZN(n17635) );
  OR2_X1 U12844 ( .A1(\pipeline/stageE/EXE_ALU/alu_shift/N202 ), .A2(
        \pipeline/EXE_controls_in_EXEcute [4]), .ZN(n17633) );
  OR2_X1 U12845 ( .A1(\pipeline/stageE/EXE_ALU/alu_shift/N202 ), .A2(
        \pipeline/EXE_controls_in_EXEcute [3]), .ZN(n17634) );
  AND2_X1 U12846 ( .A1(n14995), .A2(\pipeline/EXE_controls_in_EXEcute [6]), 
        .ZN(n17529) );
  INV_X1 U12847 ( .A(n15005), .ZN(n15001) );
  AND2_X1 U12848 ( .A1(n15165), .A2(n15166), .ZN(n17540) );
  INV_X1 U12849 ( .A(n15007), .ZN(n17551) );
  AND2_X1 U12850 ( .A1(n15145), .A2(n15138), .ZN(n17615) );
  AND3_X1 U12851 ( .A1(n17546), .A2(n15009), .A3(n15010), .ZN(n17547) );
  INV_X1 U12852 ( .A(n15161), .ZN(n15138) );
  INV_X1 U12853 ( .A(n15164), .ZN(n15165) );
  AND2_X1 U12854 ( .A1(n15011), .A2(n17533), .ZN(n17546) );
  AND2_X1 U12855 ( .A1(n15597), .A2(n15049), .ZN(n15058) );
  INV_X1 U12856 ( .A(n15445), .ZN(n15429) );
  INV_X1 U12857 ( .A(n15268), .ZN(n15281) );
  INV_X1 U12858 ( .A(n17649), .ZN(n15335) );
  INV_X1 U12859 ( .A(n15282), .ZN(n15267) );
  INV_X1 U12860 ( .A(n15015), .ZN(n17535) );
  AND3_X1 U12861 ( .A1(n17609), .A2(n17610), .A3(n17611), .ZN(n17539) );
  AND2_X1 U12862 ( .A1(\pipeline/stageE/input1_to_ALU [25]), .A2(n15234), .ZN(
        n17604) );
  AND2_X1 U12863 ( .A1(n15235), .A2(n15234), .ZN(n17605) );
  AND2_X1 U12864 ( .A1(n15235), .A2(\pipeline/stageE/input1_to_ALU [25]), .ZN(
        n17606) );
  NAND2_X1 U12865 ( .A1(n17593), .A2(n17594), .ZN(n15282) );
  INV_X1 U12866 ( .A(n17598), .ZN(n17596) );
  INV_X1 U12867 ( .A(n15314), .ZN(n15332) );
  INV_X1 U12868 ( .A(n16631), .ZN(n16630) );
  INV_X1 U12869 ( .A(n17738), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/A[16] ) );
  INV_X1 U12870 ( .A(\pipeline/stageE/input1_to_ALU [16]), .ZN(n17738) );
  AND2_X1 U12871 ( .A1(n17101), .A2(n15397), .ZN(n17592) );
  OR2_X1 U12872 ( .A1(n17101), .A2(n15397), .ZN(n17591) );
  OR2_X1 U12873 ( .A1(n15461), .A2(n15480), .ZN(n17586) );
  INV_X1 U12874 ( .A(n15461), .ZN(n17587) );
  NAND2_X1 U12875 ( .A1(n15478), .A2(n15479), .ZN(n15494) );
  OR2_X1 U12876 ( .A1(\pipeline/stageE/input1_to_ALU [7]), .A2(n15521), .ZN(
        n17583) );
  AND2_X1 U12877 ( .A1(n15525), .A2(n15540), .ZN(n17584) );
  AND3_X1 U12878 ( .A1(n17568), .A2(n17569), .A3(n17570), .ZN(
        \pipeline/stageE/input2_to_ALU[0] ) );
  NOR2_X1 U12879 ( .A1(n17387), .A2(n14982), .ZN(n17665) );
  OR2_X1 U12880 ( .A1(n17575), .A2(n17573), .ZN(
        \pipeline/stageE/EXE_ALU/alu_shift/N202 ) );
  AND2_X1 U12881 ( .A1(n16620), .A2(n13965), .ZN(n17575) );
  OR2_X1 U12882 ( .A1(n16693), .A2(\pipeline/stageE/input1_to_ALU [1]), .ZN(
        n15050) );
  AND2_X1 U12883 ( .A1(n17740), .A2(n17381), .ZN(n17576) );
  INV_X1 U12884 ( .A(n17641), .ZN(n17642) );
  INV_X1 U12885 ( .A(n16619), .ZN(n17572) );
  OR2_X1 U12886 ( .A1(n16796), .A2(n16795), .ZN(n17558) );
  INV_X1 U12887 ( .A(n16607), .ZN(n17667) );
  AND2_X1 U12888 ( .A1(\pipeline/Reg2_Addr_to_exe [3]), .A2(n17385), .ZN(
        n17549) );
  AND2_X1 U12889 ( .A1(n17314), .A2(\pipeline/Reg2_Addr_to_exe [0]), .ZN(
        n17548) );
  INV_X1 U12890 ( .A(n17346), .ZN(n17666) );
  OR2_X1 U12891 ( .A1(n14982), .A2(n17387), .ZN(n17346) );
  OR3_X1 U12892 ( .A1(n16785), .A2(n16786), .A3(n16554), .ZN(n14982) );
  INV_X1 U12893 ( .A(n17555), .ZN(n17553) );
  AND3_X1 U12894 ( .A1(n17637), .A2(n17638), .A3(n17639), .ZN(n17402) );
  INV_X1 U12895 ( .A(n14885), .ZN(n17640) );
  AND4_X1 U12896 ( .A1(n17644), .A2(n17645), .A3(n17646), .A4(n17647), .ZN(
        n16554) );
  AND2_X1 U12897 ( .A1(n17340), .A2(n17393), .ZN(n17647) );
  INV_X1 U12898 ( .A(n16585), .ZN(n16561) );
  INV_X1 U12899 ( .A(n16586), .ZN(n16805) );
  NOR2_X1 U12900 ( .A1(n16666), .A2(\pipeline/stageE/input1_to_ALU [10]), .ZN(
        n15461) );
  NOR2_X1 U12901 ( .A1(n14168), .A2(n15833), .ZN(n15610) );
  NOR2_X1 U12902 ( .A1(n15829), .A2(n15828), .ZN(n17332) );
  NOR2_X1 U12903 ( .A1(n15827), .A2(n15828), .ZN(n17330) );
  NOR2_X1 U12904 ( .A1(n15829), .A2(n15828), .ZN(n17333) );
  NOR2_X1 U12905 ( .A1(n15827), .A2(n15828), .ZN(n17331) );
  OAI21_X1 U12906 ( .B1(n17666), .B2(n17123), .A(n17327), .ZN(n16777) );
  NOR2_X1 U12907 ( .A1(n14863), .A2(n14878), .ZN(n14250) );
  NOR2_X1 U12908 ( .A1(\pipeline/EXE_controls_in_EXEcute [3]), .A2(n15584), 
        .ZN(n14964) );
  NOR2_X1 U12909 ( .A1(n16608), .A2(n17083), .ZN(n15161) );
  NOR4_X1 U12910 ( .A1(n16778), .A2(n16561), .A3(n16779), .A4(n16780), .ZN(
        n17669) );
  NOR2_X1 U12911 ( .A1(n13281), .A2(n15646), .ZN(n15611) );
  OAI21_X1 U12912 ( .B1(n16583), .B2(n16588), .A(n17703), .ZN(n13106) );
  OAI21_X1 U12913 ( .B1(n16581), .B2(n16588), .A(n17704), .ZN(n13112) );
  OAI21_X1 U12914 ( .B1(n16579), .B2(n16588), .A(n17701), .ZN(n13118) );
  OAI21_X1 U12915 ( .B1(n16576), .B2(n16588), .A(n17704), .ZN(n13124) );
  OAI21_X1 U12916 ( .B1(n16583), .B2(n16587), .A(n17703), .ZN(n13130) );
  OAI21_X1 U12917 ( .B1(n16581), .B2(n16587), .A(n17703), .ZN(n13136) );
  OAI21_X1 U12918 ( .B1(n16579), .B2(n16587), .A(n17703), .ZN(n13142) );
  OAI21_X1 U12919 ( .B1(n16576), .B2(n16587), .A(n17703), .ZN(n13148) );
  OAI21_X1 U12920 ( .B1(n16583), .B2(n16577), .A(n17705), .ZN(n13154) );
  OAI21_X1 U12921 ( .B1(n16581), .B2(n16577), .A(n17705), .ZN(n13160) );
  OAI21_X1 U12922 ( .B1(n16579), .B2(n16577), .A(n17705), .ZN(n13166) );
  OAI21_X1 U12923 ( .B1(n16576), .B2(n16577), .A(n17705), .ZN(n13172) );
  OAI21_X1 U12924 ( .B1(n16578), .B2(n16577), .A(n17705), .ZN(n13169) );
  OAI21_X1 U12925 ( .B1(n16580), .B2(n16577), .A(n17705), .ZN(n13163) );
  OAI21_X1 U12926 ( .B1(n16582), .B2(n16577), .A(n17703), .ZN(n13157) );
  NAND2_X1 U12927 ( .A1(n16584), .A2(n17643), .ZN(n16577) );
  OAI21_X1 U12928 ( .B1(n16586), .B2(n16587), .A(n17705), .ZN(n13151) );
  OAI21_X1 U12929 ( .B1(n16578), .B2(n16587), .A(n17703), .ZN(n13145) );
  OAI21_X1 U12930 ( .B1(n16580), .B2(n16587), .A(n17704), .ZN(n13139) );
  OAI21_X1 U12931 ( .B1(n16582), .B2(n16587), .A(n17703), .ZN(n13133) );
  OAI21_X1 U12932 ( .B1(n16586), .B2(n16588), .A(n17703), .ZN(n13127) );
  OAI21_X1 U12933 ( .B1(n16578), .B2(n16588), .A(n17704), .ZN(n13121) );
  OAI21_X1 U12934 ( .B1(n16580), .B2(n16588), .A(n17702), .ZN(n13115) );
  OAI21_X1 U12935 ( .B1(n16582), .B2(n16588), .A(n17704), .ZN(n13109) );
  OAI21_X1 U12936 ( .B1(n16586), .B2(n16589), .A(n17704), .ZN(n13103) );
  OAI21_X1 U12937 ( .B1(n16589), .B2(n16578), .A(n17704), .ZN(n13097) );
  NAND2_X1 U12938 ( .A1(n17703), .A2(n17650), .ZN(n13058) );
  OAI21_X1 U12939 ( .B1(n16583), .B2(n16589), .A(n17704), .ZN(n13082) );
  OAI21_X1 U12940 ( .B1(n16589), .B2(n16581), .A(n17704), .ZN(n13088) );
  NAND2_X1 U12941 ( .A1(n17703), .A2(n17651), .ZN(n13061) );
  NAND2_X1 U12942 ( .A1(n17703), .A2(n17657), .ZN(n13073) );
  NAND2_X1 U12943 ( .A1(n17703), .A2(n17661), .ZN(n13079) );
  OAI21_X1 U12944 ( .B1(n16589), .B2(n16579), .A(n17704), .ZN(n13094) );
  OAI21_X1 U12945 ( .B1(n16589), .B2(n16582), .A(n17704), .ZN(n13085) );
  NAND2_X1 U12946 ( .A1(n17703), .A2(n17658), .ZN(n13076) );
  NAND2_X1 U12947 ( .A1(n17703), .A2(n17656), .ZN(n13070) );
  OAI21_X1 U12948 ( .B1(n16589), .B2(n16576), .A(n17704), .ZN(n13100) );
  NAND2_X1 U12949 ( .A1(n17703), .A2(n17655), .ZN(n13067) );
  OAI21_X1 U12950 ( .B1(n16589), .B2(n16580), .A(n17704), .ZN(n13091) );
  NAND2_X1 U12951 ( .A1(n17703), .A2(n17654), .ZN(n13064) );
  NAND2_X1 U12952 ( .A1(n16819), .A2(n17098), .ZN(n16594) );
  NAND2_X1 U12953 ( .A1(n16822), .A2(n17098), .ZN(n16593) );
  NAND2_X1 U12954 ( .A1(n16821), .A2(n17098), .ZN(n16592) );
  NAND2_X1 U12955 ( .A1(n17660), .A2(n17098), .ZN(n16590) );
  NAND2_X1 U12956 ( .A1(n16817), .A2(n17098), .ZN(n16596) );
  NAND2_X1 U12957 ( .A1(n17125), .A2(n17098), .ZN(n16597) );
  NOR2_X1 U12958 ( .A1(n14863), .A2(n14866), .ZN(n14213) );
  NOR2_X1 U12959 ( .A1(n14864), .A2(n14867), .ZN(n14215) );
  NOR2_X1 U12960 ( .A1(n14864), .A2(n14873), .ZN(n14233) );
  NOR2_X1 U12961 ( .A1(n14865), .A2(n14873), .ZN(n14235) );
  NOR2_X1 U12962 ( .A1(n14863), .A2(n14872), .ZN(n14238) );
  NOR2_X1 U12963 ( .A1(n14863), .A2(n14873), .ZN(n14237) );
  NOR2_X1 U12964 ( .A1(n14878), .A2(n14864), .ZN(n14240) );
  NOR2_X1 U12965 ( .A1(n14865), .A2(n14878), .ZN(n14248) );
  NOR2_X1 U12966 ( .A1(n14865), .A2(n14879), .ZN(n14247) );
  NOR2_X1 U12967 ( .A1(n14879), .A2(n14863), .ZN(n14249) );
  NAND3_X1 U12968 ( .A1(n17704), .A2(n17421), .A3(
        \pipeline/EXE_controls_in_EXEcute [5]), .ZN(n14949) );
  INV_X2 U12969 ( .A(n13281), .ZN(n17705) );
  NOR3_X1 U12970 ( .A1(n15830), .A2(n15832), .A3(n15828), .ZN(n15608) );
  AOI221_X1 U12971 ( .B1(\pipeline/stageD/offset_to_jump_temp [1]), .B2(n14044), .C1(net175543), .C2(n14044), .A(n14065), .ZN(n14006) );
  NOR2_X1 U12972 ( .A1(n14862), .A2(n14863), .ZN(n17354) );
  NOR2_X1 U12973 ( .A1(n14862), .A2(n14864), .ZN(n17353) );
  NOR2_X1 U12974 ( .A1(n14860), .A2(n14867), .ZN(n17351) );
  NOR2_X1 U12975 ( .A1(n14865), .A2(n14867), .ZN(n17357) );
  NOR2_X1 U12976 ( .A1(n14862), .A2(n14863), .ZN(n17356) );
  NOR2_X1 U12977 ( .A1(n14862), .A2(n14864), .ZN(n17355) );
  NOR2_X1 U12978 ( .A1(n14860), .A2(n14867), .ZN(n17352) );
  NOR2_X1 U12979 ( .A1(n14865), .A2(n14867), .ZN(n17358) );
  NOR2_X1 U12980 ( .A1(n14862), .A2(n14863), .ZN(n17368) );
  NOR2_X1 U12981 ( .A1(n14862), .A2(n14864), .ZN(n17367) );
  AOI221_X1 U12982 ( .B1(\pipeline/stageE/EXE_ALU/alu_shift/C48/SH[1] ), .B2(
        n14968), .C1(n17741), .C2(n14981), .A(n17103), .ZN(n14975) );
  NOR2_X1 U12983 ( .A1(\pipeline/EXE_controls_in_EXEcute [2]), .A2(n15581), 
        .ZN(n17359) );
  NAND2_X1 U12984 ( .A1(\pipeline/EXE_controls_in_EXEcute [4]), .A2(n15573), 
        .ZN(n17678) );
  NOR2_X1 U12985 ( .A1(n17405), .A2(n15581), .ZN(n17360) );
  NAND2_X1 U12986 ( .A1(\pipeline/EXE_controls_in_EXEcute [4]), .A2(n15573), 
        .ZN(n17679) );
  NOR2_X1 U12987 ( .A1(n15834), .A2(n14127), .ZN(n17676) );
  NAND2_X1 U12988 ( .A1(n17674), .A2(n13944), .ZN(n17622) );
  NAND2_X1 U12989 ( .A1(\pipeline/stageF/PC_plus4/N36 ), .A2(n17108), .ZN(
        n17621) );
  AOI21_X1 U12990 ( .B1(n17631), .B2(n17632), .A(
        \pipeline/EXE_controls_in_EXEcute [6]), .ZN(n17630) );
  OAI211_X1 U12991 ( .C1(n17119), .C2(\pipeline/EXE_controls_in_EXEcute [2]), 
        .A(n17742), .B(n17633), .ZN(n17632) );
  OAI211_X1 U12992 ( .C1(n17119), .C2(
        \pipeline/stageE/EXE_ALU/add_alu/sCout[0] ), .A(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .B(n17634), .ZN(n17631) );
  NOR2_X1 U12993 ( .A1(n17405), .A2(n15581), .ZN(n17681) );
  NOR2_X1 U12994 ( .A1(\pipeline/EXE_controls_in_EXEcute [2]), .A2(n15581), 
        .ZN(n17680) );
  AOI21_X1 U12995 ( .B1(n15005), .B2(\pipeline/EXE_controls_in_EXEcute [4]), 
        .A(n17528), .ZN(n17618) );
  NOR2_X1 U12996 ( .A1(n15161), .A2(\pipeline/stageE/EXE_ALU/alu_shift/N136 ), 
        .ZN(n17608) );
  XNOR2_X1 U12997 ( .A(n17104), .B(n15137), .ZN(n17614) );
  AOI21_X1 U12998 ( .B1(n17617), .B2(n15142), .A(n15161), .ZN(n17616) );
  NAND2_X1 U12999 ( .A1(n15146), .A2(n15147), .ZN(n17617) );
  NAND2_X1 U13000 ( .A1(n15165), .A2(n15147), .ZN(n17612) );
  AOI221_X1 U13001 ( .B1(\pipeline/stageE/input1_to_ALU [19]), .B2(n15314), 
        .C1(n17649), .C2(n15316), .A(n15317), .ZN(n15296) );
  NAND2_X1 U13002 ( .A1(\pipeline/stageE/input1_to_ALU [27]), .A2(n15204), 
        .ZN(n17611) );
  NOR2_X1 U13003 ( .A1(\pipeline/stageE/input1_to_ALU [23]), .A2(n15263), .ZN(
        n17603) );
  AOI21_X1 U13004 ( .B1(n17595), .B2(n17596), .A(n17597), .ZN(n17594) );
  OAI21_X1 U13005 ( .B1(n15301), .B2(n15297), .A(n15299), .ZN(n17597) );
  NAND2_X1 U13006 ( .A1(n15319), .A2(n17599), .ZN(n17595) );
  NAND2_X1 U13007 ( .A1(n15314), .A2(\pipeline/stageE/input1_to_ALU [19]), 
        .ZN(n17599) );
  NOR2_X1 U13008 ( .A1(n17601), .A2(n17598), .ZN(n17600) );
  NAND2_X1 U13009 ( .A1(n15316), .A2(n17602), .ZN(n17598) );
  NOR2_X1 U13010 ( .A1(n15301), .A2(n15298), .ZN(n17602) );
  NAND2_X1 U13011 ( .A1(\pipeline/stageE/input1_to_ALU [11]), .A2(n15459), 
        .ZN(n17590) );
  NAND2_X1 U13012 ( .A1(\pipeline/stageE/input1_to_ALU [7]), .A2(n15521), .ZN(
        n17581) );
  NAND2_X1 U13013 ( .A1(\pipeline/EXE_controls_in_EXEcute [0]), .A2(n17400), 
        .ZN(n17570) );
  NOR2_X1 U13014 ( .A1(\pipeline/EXE_controls_in_EXEcute [0]), .A2(n13876), 
        .ZN(n17571) );
  NAND2_X1 U13015 ( .A1(n17663), .A2(\pipeline/Alu_Out_Addr_to_mem[0] ), .ZN(
        n17574) );
  NOR2_X1 U13016 ( .A1(\pipeline/EXE_controls_in_EXEcute [0]), .A2(n13848), 
        .ZN(n17577) );
  NOR2_X1 U13017 ( .A1(n17667), .A2(n17397), .ZN(n17552) );
  AOI221_X1 U13018 ( .B1(n17340), .B2(\pipeline/Reg1_Addr_to_exe [3]), .C1(
        \pipeline/regDst_to_mem[4] ), .C2(n17399), .A(n16811), .ZN(n16806) );
  NOR4_X1 U13019 ( .A1(n17559), .A2(n17560), .A3(n17561), .A4(n17562), .ZN(
        n17557) );
  OAI21_X1 U13020 ( .B1(n17385), .B2(\pipeline/Reg1_Addr_to_exe [3]), .A(
        n17563), .ZN(n17562) );
  NAND2_X1 U13021 ( .A1(n17386), .A2(\pipeline/Reg1_Addr_to_exe [4]), .ZN(
        n17563) );
  OAI21_X1 U13022 ( .B1(n17314), .B2(\pipeline/Reg1_Addr_to_exe [0]), .A(
        n17564), .ZN(n17561) );
  NAND2_X1 U13023 ( .A1(n17385), .A2(\pipeline/Reg1_Addr_to_exe [3]), .ZN(
        n17564) );
  OAI21_X1 U13024 ( .B1(\pipeline/Reg1_Addr_to_exe [1]), .B2(n17304), .A(
        n17565), .ZN(n17560) );
  NAND2_X1 U13025 ( .A1(n17314), .A2(\pipeline/Reg1_Addr_to_exe [0]), .ZN(
        n17565) );
  OAI211_X1 U13026 ( .C1(n17386), .C2(\pipeline/Reg1_Addr_to_exe [4]), .A(
        n17566), .B(n17567), .ZN(n17559) );
  NAND2_X1 U13027 ( .A1(n17304), .A2(\pipeline/Reg1_Addr_to_exe [1]), .ZN(
        n17566) );
  NAND2_X1 U13028 ( .A1(n17333), .A2(\pipeline/data_to_RF_from_WB[30] ), .ZN(
        n17639) );
  NAND2_X1 U13029 ( .A1(n17106), .A2(n17640), .ZN(n17637) );
  NOR2_X1 U13030 ( .A1(n15834), .A2(n14127), .ZN(n17675) );
  NOR2_X1 U13031 ( .A1(n16529), .A2(n16528), .ZN(n17345) );
  NOR2_X1 U13032 ( .A1(n16529), .A2(n16528), .ZN(n17337) );
  NOR2_X1 U13033 ( .A1(n16530), .A2(n16531), .ZN(n17339) );
  NOR2_X1 U13034 ( .A1(n16533), .A2(n16532), .ZN(n17335) );
  NOR2_X1 U13035 ( .A1(n16527), .A2(n16539), .ZN(n17342) );
  NOR2_X1 U13036 ( .A1(n16529), .A2(n16528), .ZN(n17336) );
  NOR2_X1 U13037 ( .A1(n16530), .A2(n16531), .ZN(n17338) );
  NOR2_X1 U13038 ( .A1(n16533), .A2(n16532), .ZN(n17334) );
  NOR2_X1 U13039 ( .A1(n16527), .A2(n16539), .ZN(n17341) );
  OAI221_X1 U13040 ( .B1(\pipeline/RegDst_to_WB[2] ), .B2(n17383), .C1(n17326), 
        .C2(\pipeline/stageD/offset_jump_sign_ext [23]), .A(n16565), .ZN(
        n16563) );
  AOI221_X1 U13041 ( .B1(\pipeline/regDst_to_mem[3] ), .B2(n17384), .C1(n17340), .C2(\pipeline/stageD/offset_jump_sign_ext [24]), .A(n16573), .ZN(n16572) );
  NOR2_X1 U13042 ( .A1(n14879), .A2(n14860), .ZN(n14245) );
  NOR2_X1 U13043 ( .A1(n14879), .A2(n14864), .ZN(n14239) );
  NOR2_X1 U13044 ( .A1(n14860), .A2(n14873), .ZN(n14227) );
  NOR2_X1 U13045 ( .A1(n14863), .A2(n14867), .ZN(n14224) );
  NOR3_X1 U13046 ( .A1(\pipeline/stageE/EXE_ALU/add_alu/sCout[0] ), .A2(
        \pipeline/EXE_controls_in_EXEcute [2]), .A3(n15586), .ZN(n14965) );
  NOR2_X1 U13047 ( .A1(n14878), .A2(n14860), .ZN(n14246) );
  NOR2_X1 U13048 ( .A1(n15348), .A2(\pipeline/stageE/input1_to_ALU [18]), .ZN(
        n16631) );
  NOR2_X1 U13049 ( .A1(n14865), .A2(n14866), .ZN(n14225) );
  NOR2_X1 U13050 ( .A1(n14864), .A2(n14866), .ZN(n14222) );
  NOR2_X1 U13051 ( .A1(n14865), .A2(n14872), .ZN(n14236) );
  NOR2_X1 U13052 ( .A1(n14864), .A2(n14872), .ZN(n14234) );
  NOR2_X1 U13053 ( .A1(n14860), .A2(n14872), .ZN(n14228) );
  NOR2_X1 U13054 ( .A1(n14865), .A2(n14862), .ZN(n14244) );
  NOR3_X1 U13055 ( .A1(\pipeline/stageE/EXE_ALU/add_alu/sCout[0] ), .A2(n17405), .A3(n15586), .ZN(n14966) );
  NOR2_X1 U13056 ( .A1(n16609), .A2(\pipeline/stageE/input1_to_ALU [29]), .ZN(
        n15164) );
  NAND2_X1 U13057 ( .A1(\pipeline/stageE/EXE_ALU/alu_shift/N202 ), .A2(n14961), 
        .ZN(n17429) );
  NAND4_X1 U13058 ( .A1(n17609), .A2(n17610), .A3(n17611), .A4(n15163), .ZN(
        n17541) );
  NAND2_X1 U13059 ( .A1(n17636), .A2(n17402), .ZN(n3989) );
  NOR2_X1 U13060 ( .A1(n17537), .A2(n17538), .ZN(n17536) );
  NAND2_X1 U13061 ( .A1(n17535), .A2(n17536), .ZN(n17534) );
  NOR3_X1 U13062 ( .A1(n15014), .A2(n15013), .A3(n17534), .ZN(n17533) );
  AOI21_X1 U13063 ( .B1(n17539), .B2(n17615), .A(n17616), .ZN(n17613) );
  XNOR2_X1 U13064 ( .A(n17539), .B(n15191), .ZN(n15011) );
  OAI21_X1 U13065 ( .B1(n17539), .B2(n15146), .A(n15145), .ZN(n15159) );
  NAND2_X1 U13066 ( .A1(n17541), .A2(n15166), .ZN(n17544) );
  NAND2_X1 U13067 ( .A1(n17541), .A2(n17540), .ZN(n17543) );
  NAND2_X1 U13068 ( .A1(n17543), .A2(n15147), .ZN(n17542) );
  XNOR2_X1 U13069 ( .A(n17544), .B(n17612), .ZN(n15010) );
  NAND3_X1 U13070 ( .A1(n15010), .A2(n15009), .A3(n17546), .ZN(n17545) );
  NAND2_X1 U13071 ( .A1(n17547), .A2(n17551), .ZN(n17619) );
  NOR2_X1 U13072 ( .A1(n17545), .A2(n17550), .ZN(n17620) );
  OAI211_X1 U13073 ( .C1(n17542), .C2(n15161), .A(n15142), .B(n13939), .ZN(
        n16598) );
  OAI22_X1 U13074 ( .A1(n17314), .A2(\pipeline/Reg2_Addr_to_exe [0]), .B1(
        n17385), .B2(\pipeline/Reg2_Addr_to_exe [3]), .ZN(n16783) );
  NOR3_X1 U13075 ( .A1(n17548), .A2(n17549), .A3(n16783), .ZN(n16782) );
  OAI221_X1 U13076 ( .B1(\pipeline/RegDst_to_WB[2] ), .B2(n17403), .C1(n17326), 
        .C2(\pipeline/Reg2_Addr_to_exe [2]), .A(n16782), .ZN(n16780) );
  NAND2_X1 U13077 ( .A1(n17411), .A2(n17551), .ZN(n17550) );
  AOI21_X1 U13078 ( .B1(n17619), .B2(n17618), .A(n17620), .ZN(n15000) );
  AOI21_X1 U13079 ( .B1(n16584), .B2(n16805), .A(n13940), .ZN(n16585) );
  AOI21_X1 U13080 ( .B1(n15123), .B2(\pipeline/data_to_RF_from_WB[1] ), .A(
        n17552), .ZN(n16699) );
  OAI22_X1 U13081 ( .A1(n17393), .A2(\pipeline/Reg2_Addr_to_exe [4]), .B1(
        n17340), .B2(\pipeline/Reg2_Addr_to_exe [3]), .ZN(n17555) );
  AOI22_X1 U13082 ( .A1(n17393), .A2(\pipeline/Reg2_Addr_to_exe [4]), .B1(
        n17340), .B2(\pipeline/Reg2_Addr_to_exe [3]), .ZN(n17554) );
  NAND2_X1 U13083 ( .A1(n17553), .A2(n17554), .ZN(n16786) );
  NOR4_X1 U13084 ( .A1(n16561), .A2(n16780), .A3(n16779), .A4(n16778), .ZN(
        n17668) );
  NOR2_X1 U13085 ( .A1(n17667), .A2(n17398), .ZN(n17556) );
  AOI21_X1 U13086 ( .B1(n17669), .B2(\pipeline/data_to_RF_from_WB[2] ), .A(
        n17556), .ZN(n16704) );
  NAND3_X1 U13087 ( .A1(n17643), .A2(n17557), .A3(n17558), .ZN(n16617) );
  XOR2_X1 U13088 ( .A(n17401), .B(\pipeline/RegDst_to_WB[2] ), .Z(n17567) );
  NAND2_X1 U13089 ( .A1(n17642), .A2(n16696), .ZN(n17568) );
  NAND2_X1 U13090 ( .A1(n16696), .A2(n17571), .ZN(n17569) );
  OAI21_X1 U13091 ( .B1(n17666), .B2(n17123), .A(n17327), .ZN(n17641) );
  OAI21_X1 U13092 ( .B1(n17105), .B2(n17396), .A(n17574), .ZN(n17573) );
  AOI21_X1 U13093 ( .B1(n17073), .B2(
        \pipeline/stageE/EXE_ALU/add_alu/sCout[0] ), .A(n17576), .ZN(n16691)
         );
  OAI22_X1 U13094 ( .A1(\pipeline/stageE/EXE_ALU/alu_shift/C48/SH[1] ), .A2(
        n17381), .B1(n17741), .B2(\pipeline/stageE/EXE_ALU/add_alu/sCout[0] ), 
        .ZN(n16693) );
  NAND2_X1 U13095 ( .A1(n15049), .A2(n15048), .ZN(n17578) );
  NAND2_X1 U13096 ( .A1(n15050), .A2(n17578), .ZN(n16690) );
  OAI21_X1 U13097 ( .B1(n15055), .B2(n16690), .A(n15053), .ZN(n16688) );
  OAI21_X1 U13098 ( .B1(n15055), .B2(n16690), .A(n15053), .ZN(n17579) );
  NAND2_X1 U13099 ( .A1(n15566), .A2(n15569), .ZN(n16682) );
  NAND2_X1 U13100 ( .A1(n16682), .A2(n15568), .ZN(n15541) );
  NAND3_X1 U13101 ( .A1(n17582), .A2(n15527), .A3(n17583), .ZN(n17580) );
  OAI21_X1 U13102 ( .B1(n15541), .B2(n15542), .A(n17584), .ZN(n17582) );
  NAND2_X1 U13103 ( .A1(n17580), .A2(n17581), .ZN(n15508) );
  NAND2_X1 U13104 ( .A1(n15508), .A2(n15509), .ZN(n15478) );
  NAND3_X1 U13105 ( .A1(n17585), .A2(n15463), .A3(n17586), .ZN(n16664) );
  NAND3_X1 U13106 ( .A1(n15494), .A2(n15495), .A3(n17587), .ZN(n17585) );
  NAND2_X1 U13107 ( .A1(n16664), .A2(\pipeline/stageE/input1_to_ALU [11]), 
        .ZN(n17588) );
  NAND2_X1 U13108 ( .A1(n16664), .A2(n15459), .ZN(n17589) );
  NAND3_X1 U13109 ( .A1(n15367), .A2(n15383), .A3(n16630), .ZN(n17601) );
  NAND2_X1 U13110 ( .A1(n15368), .A2(n17600), .ZN(n17593) );
  OAI221_X1 U13111 ( .B1(n15248), .B2(n17117), .C1(n15248), .C2(n16613), .A(
        n15250), .ZN(n15235) );
  XOR2_X1 U13112 ( .A(n17078), .B(n15204), .Z(n17607) );
  XNOR2_X1 U13113 ( .A(n15205), .B(n17607), .ZN(n15014) );
  NAND2_X1 U13114 ( .A1(n15205), .A2(\pipeline/stageE/input1_to_ALU [27]), 
        .ZN(n17609) );
  NAND2_X1 U13115 ( .A1(n15205), .A2(n15204), .ZN(n17610) );
  XNOR2_X1 U13116 ( .A(n17613), .B(n17614), .ZN(n15007) );
  OAI211_X1 U13117 ( .C1(n15046), .C2(n14949), .A(n17429), .B(n17629), .ZN(
        n17628) );
  AOI21_X1 U13118 ( .B1(\pipeline/stageE/EXE_ALU/alu_shift/N234 ), .B2(n17681), 
        .A(n17628), .ZN(n17627) );
  NAND2_X1 U13119 ( .A1(\pipeline/stageE/EXE_ALU/alu_shift/N39 ), .A2(n17149), 
        .ZN(n17626) );
  NAND2_X1 U13120 ( .A1(n17624), .A2(n17635), .ZN(n17623) );
  NAND2_X1 U13121 ( .A1(n17630), .A2(n14995), .ZN(n17629) );
  NAND2_X1 U13122 ( .A1(\pipeline/stageE/EXE_ALU/alu_shift/N7 ), .A2(n14965), 
        .ZN(n17625) );
  NAND2_X1 U13123 ( .A1(\pipeline/stageE/EXE_ALU/alu_shift/N137 ), .A2(n17680), 
        .ZN(n17624) );
  NAND2_X1 U13124 ( .A1(\pipeline/stageD/target_Jump_temp [30]), .A2(n17675), 
        .ZN(n17636) );
  OAI221_X1 U13125 ( .B1(\pipeline/stageD/offset_to_jump_temp [7]), .B2(
        \pipeline/stageD/offset_to_jump_temp [2]), .C1(
        \pipeline/stageD/offset_to_jump_temp [7]), .C2(n17406), .A(
        \pipeline/cu_pipeline/N89 ), .ZN(n14072) );
  NOR4_X1 U13126 ( .A1(\pipeline/stageD/offset_to_jump_temp [3]), .A2(
        \pipeline/stageD/offset_to_jump_temp [4]), .A3(
        \pipeline/stageD/offset_to_jump_temp [2]), .A4(n17350), .ZN(n13990) );
  AOI22_X1 U13127 ( .A1(n17671), .A2(\pipeline/stageD/offset_to_jump_temp [2]), 
        .B1(n17107), .B2(InstrFetched[2]), .ZN(n15623) );
  NAND4_X1 U13128 ( .A1(\pipeline/stageD/offset_to_jump_temp [3]), .A2(
        \pipeline/stageD/offset_to_jump_temp [5]), .A3(
        \pipeline/stageD/offset_to_jump_temp [2]), .A4(n17406), .ZN(n14180) );
  NOR3_X1 U13129 ( .A1(\pipeline/stageD/offset_to_jump_temp [2]), .A2(n17410), 
        .A3(n17350), .ZN(n14179) );
  AOI22_X1 U13130 ( .A1(n17671), .A2(\pipeline/nextPC_IFID_DEC[0] ), .B1(
        n17673), .B2(\pipeline/stageF/PC_plus4/N7 ), .ZN(n15773) );
  AOI22_X1 U13131 ( .A1(n17663), .A2(\pipeline/Alu_Out_Addr_to_mem[29] ), .B1(
        n16620), .B2(n13956), .ZN(n16770) );
  AOI22_X1 U13132 ( .A1(n17663), .A2(\pipeline/Alu_Out_Addr_to_mem[28] ), .B1(
        n16620), .B2(n13962), .ZN(n16766) );
  AOI22_X1 U13133 ( .A1(n17663), .A2(\pipeline/Alu_Out_Addr_to_mem[23] ), .B1(
        n16620), .B2(n13952), .ZN(n16753) );
  AOI22_X1 U13134 ( .A1(n17663), .A2(\pipeline/Alu_Out_Addr_to_mem[19] ), .B1(
        n16620), .B2(n13948), .ZN(n16637) );
  AOI22_X1 U13135 ( .A1(n17663), .A2(\pipeline/Alu_Out_Addr_to_mem[15] ), .B1(
        n16620), .B2(n13959), .ZN(n16733) );
  AOI22_X1 U13136 ( .A1(n17663), .A2(\pipeline/Alu_Out_Addr_to_mem[18] ), .B1(
        n16620), .B2(n13947), .ZN(n16734) );
  AOI22_X1 U13137 ( .A1(n17663), .A2(\pipeline/Alu_Out_Addr_to_mem[16] ), .B1(
        n16620), .B2(n13804), .ZN(n16641) );
  AOI22_X1 U13138 ( .A1(n17663), .A2(\pipeline/Alu_Out_Addr_to_mem[9] ), .B1(
        n16620), .B2(n13820), .ZN(n16671) );
  AOI22_X1 U13139 ( .A1(n17663), .A2(\pipeline/Alu_Out_Addr_to_mem[8] ), .B1(
        n16620), .B2(n13964), .ZN(n16720) );
  AOI22_X1 U13140 ( .A1(n17663), .A2(\pipeline/Alu_Out_Addr_to_mem[1] ), .B1(
        n16620), .B2(n13847), .ZN(n16701) );
  XNOR2_X1 U13141 ( .A(\pipeline/stageE/EXE_ALU/add_alu/sCout[0] ), .B(n15133), 
        .ZN(n15137) );
  XNOR2_X1 U13142 ( .A(n15493), .B(n15494), .ZN(n15035) );
  OAI221_X1 U13143 ( .B1(n15477), .B2(n15478), .C1(n15477), .C2(n15479), .A(
        n15480), .ZN(n15476) );
  AOI22_X1 U13144 ( .A1(n17665), .A2(\pipeline/Alu_Out_Addr_to_mem[29] ), .B1(
        n17123), .B2(\pipeline/data_to_RF_from_WB[29] ), .ZN(n16773) );
  AOI22_X1 U13145 ( .A1(n17666), .A2(\pipeline/Alu_Out_Addr_to_mem[25] ), .B1(
        n17123), .B2(\pipeline/data_to_RF_from_WB[25] ), .ZN(n16757) );
  AOI22_X1 U13146 ( .A1(n17666), .A2(\pipeline/Alu_Out_Addr_to_mem[23] ), .B1(
        n17123), .B2(\pipeline/data_to_RF_from_WB[23] ), .ZN(n16752) );
  AOI22_X1 U13147 ( .A1(n17666), .A2(\pipeline/Alu_Out_Addr_to_mem[16] ), .B1(
        n17123), .B2(\pipeline/data_to_RF_from_WB[16] ), .ZN(n16640) );
  AOI22_X1 U13148 ( .A1(n17665), .A2(\pipeline/Alu_Out_Addr_to_mem[12] ), .B1(
        n17123), .B2(\pipeline/data_to_RF_from_WB[12] ), .ZN(n16663) );
  NOR2_X1 U13149 ( .A1(n17340), .A2(n14129), .ZN(\pipeline/MEMWB_Stage/N46 )
         );
  OAI22_X1 U13150 ( .A1(n17304), .A2(
        \pipeline/stageD/offset_jump_sign_ext [22]), .B1(n17386), .B2(
        \pipeline/stageD/offset_jump_sign_ext [31]), .ZN(n16568) );
  AOI22_X1 U13151 ( .A1(n17304), .A2(\pipeline/Reg2_Addr_to_exe [1]), .B1(
        \pipeline/Reg2_Addr_to_exe [4]), .B2(n17386), .ZN(n16784) );
  NAND3_X1 U13152 ( .A1(n15368), .A2(n15367), .A3(n15383), .ZN(n17648) );
  AOI22_X1 U13153 ( .A1(\pipeline/data_to_RF_from_WB[0] ), .A2(n17123), .B1(
        \pipeline/Alu_Out_Addr_to_mem[0] ), .B2(n17665), .ZN(n16696) );
  OAI21_X1 U13154 ( .B1(n15596), .B2(\pipeline/stageE/EXE_ALU/alu_shift/N202 ), 
        .A(n15050), .ZN(n15597) );
  NOR2_X1 U13155 ( .A1(n16631), .A2(n17648), .ZN(n17649) );
  NAND2_X1 U13156 ( .A1(n15049), .A2(n15050), .ZN(n15047) );
  NAND2_X1 U13157 ( .A1(n16806), .A2(n16807), .ZN(n16796) );
  NAND2_X1 U13158 ( .A1(n15049), .A2(n15595), .ZN(n15056) );
  NOR4_X1 U13159 ( .A1(n16778), .A2(n16561), .A3(n16779), .A4(n16780), .ZN(
        n15123) );
  XNOR2_X1 U13160 ( .A(n15554), .B(n15541), .ZN(n15042) );
  AOI21_X1 U13161 ( .B1(n15540), .B2(n15541), .A(n15542), .ZN(n15526) );
  NOR2_X1 U13162 ( .A1(n16554), .A2(n16555), .ZN(n14103) );
  OAI221_X1 U13163 ( .B1(\pipeline/regDst_to_mem[4] ), .B2(n17328), .C1(n17393), .C2(\pipeline/stageD/offset_jump_sign_ext [31]), .A(n16574), .ZN(n16573) );
  OAI22_X1 U13164 ( .A1(n17340), .A2(\pipeline/Reg1_Addr_to_exe [3]), .B1(
        n17399), .B2(\pipeline/regDst_to_mem[4] ), .ZN(n16811) );
  OAI22_X1 U13165 ( .A1(\pipeline/stageE/EXE_ALU/alu_shift/N202 ), .A2(
        \pipeline/stageE/EXE_ALU/alu_shift/C48/SH[0] ), .B1(n17742), .B2(
        n17119), .ZN(n15046) );
  AOI22_X1 U13166 ( .A1(\pipeline/stageE/EXE_ALU/add_alu/sCout[0] ), .A2(
        \pipeline/stageE/input2_to_ALU[0] ), .B1(n17742), .B2(n17381), .ZN(
        n15596) );
  AOI21_X1 U13167 ( .B1(n15416), .B2(n16652), .A(n15413), .ZN(n16650) );
  OAI211_X1 U13168 ( .C1(net175543), .C2(n13990), .A(
        \pipeline/stageD/offset_to_jump_temp [1]), .B(
        \pipeline/cu_pipeline/N89 ), .ZN(n14071) );
  AOI22_X1 U13169 ( .A1(n17671), .A2(net175543), .B1(n15601), .B2(
        InstrFetched[0]), .ZN(n15621) );
  NOR2_X1 U13170 ( .A1(net175543), .A2(n17406), .ZN(n14051) );
  NOR2_X1 U13171 ( .A1(\pipeline/stageD/offset_to_jump_temp [1]), .A2(
        net175543), .ZN(n14032) );
  XNOR2_X1 U13172 ( .A(n15047), .B(n15048), .ZN(n14970) );
  NOR3_X1 U13173 ( .A1(\pipeline/stageE/EXE_ALU/alu_shift/C48/SH[1] ), .A2(
        \pipeline/stageE/input1_to_ALU [1]), .A3(n17678), .ZN(n14974) );
  AOI211_X1 U13174 ( .C1(n14993), .C2(n15007), .A(n15126), .B(n15127), .ZN(
        n15125) );
  XNOR2_X1 U13175 ( .A(n15217), .B(n15218), .ZN(n15015) );
  XNOR2_X1 U13176 ( .A(n15234), .B(n15235), .ZN(n15233) );
  NAND2_X1 U13177 ( .A1(n15445), .A2(n15446), .ZN(n16657) );
  NOR2_X1 U13178 ( .A1(n16650), .A2(n15398), .ZN(n16646) );
endmodule

