
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_DLX;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity DLX is

   port( Clk, Rst : in std_logic;  exception : out std_logic);

end DLX;

architecture SYN_struct of DLX is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X2
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X2
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X2
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   component IRAM
      port( ck, Rst : in std_logic;  Addr : in std_logic_vector (31 downto 0); 
            Dout : out std_logic_vector (31 downto 0));
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component TINV_X1
      port( I, EN : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal addr_to_iram_31_port, addr_to_iram_30_port, addr_to_iram_29_port, 
      addr_to_iram_28_port, addr_to_iram_27_port, addr_to_iram_26_port, 
      addr_to_iram_25_port, addr_to_iram_24_port, addr_to_iram_23_port, 
      addr_to_iram_22_port, addr_to_iram_21_port, addr_to_iram_20_port, 
      addr_to_iram_19_port, addr_to_iram_18_port, addr_to_iram_17_port, 
      addr_to_iram_16_port, addr_to_iram_15_port, addr_to_iram_14_port, 
      addr_to_iram_13_port, addr_to_iram_12_port, addr_to_iram_11_port, 
      addr_to_iram_10_port, addr_to_iram_9_port, addr_to_iram_8_port, 
      addr_to_iram_7_port, addr_to_iram_6_port, addr_to_iram_5_port, 
      addr_to_iram_4_port, addr_to_iram_3_port, addr_to_iram_2_port, 
      InstrFetched_31_port, InstrFetched_30_port, InstrFetched_29_port, 
      InstrFetched_28_port, InstrFetched_27_port, InstrFetched_26_port, 
      InstrFetched_25_port, InstrFetched_24_port, InstrFetched_23_port, 
      InstrFetched_22_port, InstrFetched_21_port, InstrFetched_20_port, 
      InstrFetched_19_port, InstrFetched_18_port, InstrFetched_17_port, 
      InstrFetched_16_port, InstrFetched_15_port, InstrFetched_14_port, 
      InstrFetched_13_port, InstrFetched_12_port, InstrFetched_11_port, 
      InstrFetched_10_port, InstrFetched_9_port, InstrFetched_8_port, 
      InstrFetched_7_port, InstrFetched_6_port, InstrFetched_5_port, 
      InstrFetched_4_port, InstrFetched_3_port, InstrFetched_2_port, 
      InstrFetched_1_port, InstrFetched_0_port, data_from_dram_31_port, 
      data_from_dram_30_port, data_from_dram_29_port, data_from_dram_28_port, 
      data_from_dram_27_port, data_from_dram_26_port, data_from_dram_25_port, 
      data_from_dram_24_port, data_from_dram_23_port, data_from_dram_22_port, 
      data_from_dram_21_port, data_from_dram_20_port, data_from_dram_19_port, 
      data_from_dram_18_port, data_from_dram_17_port, data_from_dram_16_port, 
      data_from_dram_15_port, data_from_dram_14_port, data_from_dram_13_port, 
      data_from_dram_12_port, data_from_dram_11_port, data_from_dram_10_port, 
      data_from_dram_9_port, data_from_dram_8_port, data_from_dram_7_port, 
      data_from_dram_6_port, data_from_dram_5_port, data_from_dram_4_port, 
      data_from_dram_3_port, data_from_dram_2_port, data_from_dram_1_port, 
      data_from_dram_0_port, read_notWrite, addr_to_dataRam_4_port, 
      addr_to_dataRam_3_port, addr_to_dataRam_2_port, pipeline_Forward_sw1_mux,
      pipeline_regDst_to_mem_0_port, pipeline_regDst_to_mem_1_port, 
      pipeline_regDst_to_mem_3_port, pipeline_regDst_to_mem_4_port, 
      pipeline_MEM_controls_in_MEM_1_port, pipeline_WB_controls_in_MEMWB_0_port
      , pipeline_WB_controls_in_MEMWB_1_port, pipeline_immediate_to_exe_1_port,
      pipeline_immediate_to_exe_2_port, pipeline_immediate_to_exe_3_port, 
      pipeline_immediate_to_exe_4_port, pipeline_immediate_to_exe_5_port, 
      pipeline_immediate_to_exe_6_port, pipeline_immediate_to_exe_7_port, 
      pipeline_immediate_to_exe_8_port, pipeline_immediate_to_exe_9_port, 
      pipeline_immediate_to_exe_10_port, pipeline_immediate_to_exe_11_port, 
      pipeline_immediate_to_exe_12_port, pipeline_immediate_to_exe_13_port, 
      pipeline_immediate_to_exe_14_port, pipeline_immediate_to_exe_15_port, 
      pipeline_immediate_to_exe_16_port, pipeline_immediate_to_exe_17_port, 
      pipeline_immediate_to_exe_18_port, pipeline_immediate_to_exe_19_port, 
      pipeline_immediate_to_exe_20_port, pipeline_immediate_to_exe_21_port, 
      pipeline_immediate_to_exe_22_port, pipeline_immediate_to_exe_23_port, 
      pipeline_immediate_to_exe_24_port, pipeline_immediate_to_exe_25_port, 
      pipeline_immediate_to_exe_26_port, pipeline_immediate_to_exe_27_port, 
      pipeline_immediate_to_exe_28_port, pipeline_immediate_to_exe_29_port, 
      pipeline_immediate_to_exe_30_port, pipeline_immediate_to_exe_31_port, 
      pipeline_Reg2_Addr_to_exe_0_port, pipeline_Reg2_Addr_to_exe_1_port, 
      pipeline_Reg2_Addr_to_exe_2_port, pipeline_Reg2_Addr_to_exe_3_port, 
      pipeline_Reg2_Addr_to_exe_4_port, pipeline_Reg1_Addr_to_exe_0_port, 
      pipeline_Reg1_Addr_to_exe_1_port, pipeline_Reg1_Addr_to_exe_2_port, 
      pipeline_Reg1_Addr_to_exe_3_port, pipeline_Reg1_Addr_to_exe_4_port, 
      pipeline_EXE_controls_in_EXEcute_0_port, 
      pipeline_EXE_controls_in_EXEcute_2_port, 
      pipeline_EXE_controls_in_EXEcute_3_port, 
      pipeline_EXE_controls_in_EXEcute_4_port, 
      pipeline_EXE_controls_in_EXEcute_5_port, 
      pipeline_EXE_controls_in_EXEcute_6_port, 
      pipeline_EXE_controls_in_EXEcute_7_port, 
      pipeline_MEM_controls_in_EXMEM_1_port, 
      pipeline_WB_controls_in_EXMEM_1_port, pipeline_WB_controls_in_IDEX_0_port
      , pipeline_RegDst_to_WB_0_port, pipeline_RegDst_to_WB_1_port, 
      pipeline_RegDst_to_WB_2_port, pipeline_RegDst_to_WB_3_port, 
      pipeline_RegDst_to_WB_4_port, pipeline_EXE_controls_in_IDEX_0_port, 
      pipeline_EXE_controls_in_IDEX_1_port, 
      pipeline_EXE_controls_in_IDEX_2_port, 
      pipeline_EXE_controls_in_IDEX_3_port, 
      pipeline_EXE_controls_in_IDEX_4_port, 
      pipeline_EXE_controls_in_IDEX_5_port, 
      pipeline_EXE_controls_in_IDEX_6_port, 
      pipeline_EXE_controls_in_IDEX_7_port, 
      pipeline_EXE_controls_in_IDEX_8_port, pipeline_data_to_RF_from_WB_0_port,
      pipeline_data_to_RF_from_WB_1_port, pipeline_data_to_RF_from_WB_2_port, 
      pipeline_data_to_RF_from_WB_3_port, pipeline_data_to_RF_from_WB_4_port, 
      pipeline_data_to_RF_from_WB_5_port, pipeline_data_to_RF_from_WB_6_port, 
      pipeline_data_to_RF_from_WB_7_port, pipeline_data_to_RF_from_WB_8_port, 
      pipeline_data_to_RF_from_WB_9_port, pipeline_data_to_RF_from_WB_10_port, 
      pipeline_data_to_RF_from_WB_11_port, pipeline_data_to_RF_from_WB_12_port,
      pipeline_data_to_RF_from_WB_13_port, pipeline_data_to_RF_from_WB_14_port,
      pipeline_data_to_RF_from_WB_15_port, pipeline_data_to_RF_from_WB_16_port,
      pipeline_data_to_RF_from_WB_17_port, pipeline_data_to_RF_from_WB_18_port,
      pipeline_data_to_RF_from_WB_19_port, pipeline_data_to_RF_from_WB_20_port,
      pipeline_data_to_RF_from_WB_21_port, pipeline_data_to_RF_from_WB_22_port,
      pipeline_data_to_RF_from_WB_23_port, pipeline_data_to_RF_from_WB_24_port,
      pipeline_data_to_RF_from_WB_25_port, pipeline_data_to_RF_from_WB_26_port,
      pipeline_data_to_RF_from_WB_27_port, pipeline_data_to_RF_from_WB_28_port,
      pipeline_data_to_RF_from_WB_29_port, pipeline_data_to_RF_from_WB_30_port,
      pipeline_data_to_RF_from_WB_31_port, pipeline_Alu_Out_Addr_to_mem_0_port,
      pipeline_Alu_Out_Addr_to_mem_1_port, pipeline_Alu_Out_Addr_to_mem_2_port,
      pipeline_Alu_Out_Addr_to_mem_3_port, pipeline_Alu_Out_Addr_to_mem_4_port,
      pipeline_Alu_Out_Addr_to_mem_5_port, pipeline_Alu_Out_Addr_to_mem_6_port,
      pipeline_Alu_Out_Addr_to_mem_7_port, pipeline_Alu_Out_Addr_to_mem_8_port,
      pipeline_Alu_Out_Addr_to_mem_9_port, pipeline_Alu_Out_Addr_to_mem_10_port
      , pipeline_Alu_Out_Addr_to_mem_11_port, 
      pipeline_Alu_Out_Addr_to_mem_12_port, 
      pipeline_Alu_Out_Addr_to_mem_13_port, 
      pipeline_Alu_Out_Addr_to_mem_14_port, 
      pipeline_Alu_Out_Addr_to_mem_15_port, 
      pipeline_Alu_Out_Addr_to_mem_16_port, 
      pipeline_Alu_Out_Addr_to_mem_17_port, 
      pipeline_Alu_Out_Addr_to_mem_18_port, 
      pipeline_Alu_Out_Addr_to_mem_19_port, 
      pipeline_Alu_Out_Addr_to_mem_20_port, 
      pipeline_Alu_Out_Addr_to_mem_21_port, 
      pipeline_Alu_Out_Addr_to_mem_22_port, 
      pipeline_Alu_Out_Addr_to_mem_23_port, 
      pipeline_Alu_Out_Addr_to_mem_24_port, 
      pipeline_Alu_Out_Addr_to_mem_25_port, 
      pipeline_Alu_Out_Addr_to_mem_26_port, 
      pipeline_Alu_Out_Addr_to_mem_27_port, 
      pipeline_Alu_Out_Addr_to_mem_28_port, 
      pipeline_Alu_Out_Addr_to_mem_29_port, 
      pipeline_Alu_Out_Addr_to_mem_30_port, 
      pipeline_Alu_Out_Addr_to_mem_31_port, pipeline_inst_IFID_DEC_26_port, 
      pipeline_inst_IFID_DEC_27_port, pipeline_inst_IFID_DEC_28_port, 
      pipeline_inst_IFID_DEC_29_port, pipeline_inst_IFID_DEC_30_port, 
      pipeline_inst_IFID_DEC_31_port, pipeline_nextPC_IFID_DEC_0_port, 
      pipeline_nextPC_IFID_DEC_1_port, pipeline_nextPC_IFID_DEC_2_port, 
      pipeline_nextPC_IFID_DEC_3_port, pipeline_nextPC_IFID_DEC_4_port, 
      pipeline_nextPC_IFID_DEC_5_port, pipeline_nextPC_IFID_DEC_6_port, 
      pipeline_nextPC_IFID_DEC_7_port, pipeline_nextPC_IFID_DEC_8_port, 
      pipeline_nextPC_IFID_DEC_9_port, pipeline_nextPC_IFID_DEC_10_port, 
      pipeline_nextPC_IFID_DEC_11_port, pipeline_nextPC_IFID_DEC_12_port, 
      pipeline_nextPC_IFID_DEC_13_port, pipeline_nextPC_IFID_DEC_14_port, 
      pipeline_nextPC_IFID_DEC_15_port, pipeline_nextPC_IFID_DEC_16_port, 
      pipeline_nextPC_IFID_DEC_17_port, pipeline_nextPC_IFID_DEC_18_port, 
      pipeline_nextPC_IFID_DEC_19_port, pipeline_nextPC_IFID_DEC_20_port, 
      pipeline_nextPC_IFID_DEC_21_port, pipeline_nextPC_IFID_DEC_22_port, 
      pipeline_nextPC_IFID_DEC_23_port, pipeline_nextPC_IFID_DEC_24_port, 
      pipeline_nextPC_IFID_DEC_25_port, pipeline_nextPC_IFID_DEC_26_port, 
      pipeline_nextPC_IFID_DEC_27_port, pipeline_nextPC_IFID_DEC_28_port, 
      pipeline_nextPC_IFID_DEC_29_port, pipeline_nextPC_IFID_DEC_30_port, 
      pipeline_stall, pipeline_stageF_PC_plus4_N37, 
      pipeline_stageF_PC_plus4_N36, pipeline_stageF_PC_plus4_N35, 
      pipeline_stageF_PC_plus4_N34, pipeline_stageF_PC_plus4_N33, 
      pipeline_stageF_PC_plus4_N32, pipeline_stageF_PC_plus4_N31, 
      pipeline_stageF_PC_plus4_N30, pipeline_stageF_PC_plus4_N29, 
      pipeline_stageF_PC_plus4_N28, pipeline_stageF_PC_plus4_N27, 
      pipeline_stageF_PC_plus4_N26, pipeline_stageF_PC_plus4_N25, 
      pipeline_stageF_PC_plus4_N24, pipeline_stageF_PC_plus4_N23, 
      pipeline_stageF_PC_plus4_N22, pipeline_stageF_PC_plus4_N21, 
      pipeline_stageF_PC_plus4_N20, pipeline_stageF_PC_plus4_N19, 
      pipeline_stageF_PC_plus4_N18, pipeline_stageF_PC_plus4_N17, 
      pipeline_stageF_PC_plus4_N16, pipeline_stageF_PC_plus4_N15, 
      pipeline_stageF_PC_plus4_N14, pipeline_stageF_PC_plus4_N13, 
      pipeline_stageF_PC_plus4_N12, pipeline_stageF_PC_plus4_N11, 
      pipeline_stageF_PC_plus4_N10, pipeline_stageF_PC_plus4_N9, 
      pipeline_stageF_PC_plus4_N8, pipeline_stageF_PC_plus4_N7, 
      pipeline_stageF_PC_reg_N31, pipeline_stageF_PC_reg_N30, 
      pipeline_stageF_PC_reg_N29, pipeline_stageF_PC_reg_N28, 
      pipeline_stageF_PC_reg_N27, pipeline_stageF_PC_reg_N26, 
      pipeline_stageF_PC_reg_N25, pipeline_stageF_PC_reg_N24, 
      pipeline_stageF_PC_reg_N23, pipeline_stageF_PC_reg_N22, 
      pipeline_stageF_PC_reg_N21, pipeline_stageF_PC_reg_N20, 
      pipeline_stageF_PC_reg_N19, pipeline_stageF_PC_reg_N18, 
      pipeline_stageF_PC_reg_N17, pipeline_stageF_PC_reg_N16, 
      pipeline_stageF_PC_reg_N15, pipeline_stageF_PC_reg_N14, 
      pipeline_stageF_PC_reg_N13, pipeline_stageF_PC_reg_N12, 
      pipeline_stageF_PC_reg_N11, pipeline_stageF_PC_reg_N10, 
      pipeline_stageF_PC_reg_N9, pipeline_stageF_PC_reg_N8, 
      pipeline_stageF_PC_reg_N7, pipeline_stageF_PC_reg_N6, 
      pipeline_stageF_PC_reg_N5, pipeline_stageF_PC_reg_N4, 
      pipeline_stageF_PC_reg_N3, pipeline_stageF_PC_reg_N2, 
      pipeline_stageF_PC_reg_N1, pipeline_stageF_PC_reg_N0, 
      pipeline_stageD_target_Jump_temp_0_port, 
      pipeline_stageD_target_Jump_temp_1_port, 
      pipeline_stageD_target_Jump_temp_2_port, 
      pipeline_stageD_target_Jump_temp_3_port, 
      pipeline_stageD_target_Jump_temp_4_port, 
      pipeline_stageD_target_Jump_temp_5_port, 
      pipeline_stageD_target_Jump_temp_6_port, 
      pipeline_stageD_target_Jump_temp_7_port, 
      pipeline_stageD_target_Jump_temp_8_port, 
      pipeline_stageD_target_Jump_temp_9_port, 
      pipeline_stageD_target_Jump_temp_10_port, 
      pipeline_stageD_target_Jump_temp_11_port, 
      pipeline_stageD_target_Jump_temp_12_port, 
      pipeline_stageD_target_Jump_temp_13_port, 
      pipeline_stageD_target_Jump_temp_14_port, 
      pipeline_stageD_target_Jump_temp_15_port, 
      pipeline_stageD_target_Jump_temp_16_port, 
      pipeline_stageD_target_Jump_temp_17_port, 
      pipeline_stageD_target_Jump_temp_18_port, 
      pipeline_stageD_target_Jump_temp_19_port, 
      pipeline_stageD_target_Jump_temp_20_port, 
      pipeline_stageD_target_Jump_temp_21_port, 
      pipeline_stageD_target_Jump_temp_22_port, 
      pipeline_stageD_target_Jump_temp_23_port, 
      pipeline_stageD_target_Jump_temp_24_port, 
      pipeline_stageD_target_Jump_temp_25_port, 
      pipeline_stageD_target_Jump_temp_26_port, 
      pipeline_stageD_target_Jump_temp_27_port, 
      pipeline_stageD_target_Jump_temp_28_port, 
      pipeline_stageD_target_Jump_temp_29_port, 
      pipeline_stageD_target_Jump_temp_30_port, 
      pipeline_stageD_target_Jump_temp_31_port, 
      pipeline_stageD_offset_to_jump_temp_1_port, 
      pipeline_stageD_offset_to_jump_temp_2_port, 
      pipeline_stageD_offset_to_jump_temp_3_port, 
      pipeline_stageD_offset_to_jump_temp_4_port, 
      pipeline_stageD_offset_to_jump_temp_5_port, 
      pipeline_stageD_offset_to_jump_temp_6_port, 
      pipeline_stageD_offset_to_jump_temp_7_port, 
      pipeline_stageD_offset_to_jump_temp_8_port, 
      pipeline_stageD_offset_to_jump_temp_9_port, 
      pipeline_stageD_offset_to_jump_temp_10_port, 
      pipeline_stageD_offset_to_jump_temp_11_port, 
      pipeline_stageD_offset_to_jump_temp_12_port, 
      pipeline_stageD_offset_to_jump_temp_13_port, 
      pipeline_stageD_offset_to_jump_temp_14_port, 
      pipeline_stageD_offset_to_jump_temp_15_port, 
      pipeline_stageD_offset_to_jump_temp_16_port, 
      pipeline_stageD_offset_to_jump_temp_17_port, 
      pipeline_stageD_offset_to_jump_temp_18_port, 
      pipeline_stageD_offset_to_jump_temp_19_port, 
      pipeline_stageD_offset_to_jump_temp_20_port, 
      pipeline_stageD_offset_to_jump_temp_21_port, 
      pipeline_stageD_offset_to_jump_temp_22_port, 
      pipeline_stageD_offset_to_jump_temp_23_port, 
      pipeline_stageD_offset_to_jump_temp_24_port, 
      pipeline_stageD_offset_to_jump_temp_30_port, 
      pipeline_stageD_offset_jump_sign_ext_16_port, 
      pipeline_stageD_offset_jump_sign_ext_17_port, 
      pipeline_stageD_offset_jump_sign_ext_18_port, 
      pipeline_stageD_offset_jump_sign_ext_19_port, 
      pipeline_stageD_offset_jump_sign_ext_20_port, 
      pipeline_stageD_offset_jump_sign_ext_21_port, 
      pipeline_stageD_offset_jump_sign_ext_22_port, 
      pipeline_stageD_offset_jump_sign_ext_23_port, 
      pipeline_stageD_offset_jump_sign_ext_24_port, 
      pipeline_stageD_offset_jump_sign_ext_31_port, 
      pipeline_stageD_evaluate_jump_target_N63, 
      pipeline_stageD_evaluate_jump_target_N62, 
      pipeline_stageD_evaluate_jump_target_N61, 
      pipeline_stageD_evaluate_jump_target_N60, 
      pipeline_stageD_evaluate_jump_target_N59, 
      pipeline_stageD_evaluate_jump_target_N58, 
      pipeline_stageD_evaluate_jump_target_N57, 
      pipeline_stageD_evaluate_jump_target_N56, 
      pipeline_stageD_evaluate_jump_target_N55, 
      pipeline_stageD_evaluate_jump_target_N54, 
      pipeline_stageD_evaluate_jump_target_N53, 
      pipeline_stageD_evaluate_jump_target_N52, 
      pipeline_stageD_evaluate_jump_target_N51, 
      pipeline_stageD_evaluate_jump_target_N50, 
      pipeline_stageD_evaluate_jump_target_N49, 
      pipeline_stageD_evaluate_jump_target_N48, 
      pipeline_stageD_evaluate_jump_target_N47, 
      pipeline_stageD_evaluate_jump_target_N46, 
      pipeline_stageD_evaluate_jump_target_N45, 
      pipeline_stageD_evaluate_jump_target_N44, 
      pipeline_stageD_evaluate_jump_target_N43, 
      pipeline_stageD_evaluate_jump_target_N42, 
      pipeline_stageD_evaluate_jump_target_N41, 
      pipeline_stageD_evaluate_jump_target_N40, 
      pipeline_stageD_evaluate_jump_target_N39, 
      pipeline_stageD_evaluate_jump_target_N38, 
      pipeline_stageD_evaluate_jump_target_N37, 
      pipeline_stageD_evaluate_jump_target_N36, 
      pipeline_stageD_evaluate_jump_target_N35, 
      pipeline_stageD_evaluate_jump_target_N34, 
      pipeline_stageD_evaluate_jump_target_N33, 
      pipeline_RegFile_DEC_WB_RegBank_31_0_port, 
      pipeline_RegFile_DEC_WB_RegBank_31_1_port, 
      pipeline_RegFile_DEC_WB_RegBank_31_2_port, 
      pipeline_RegFile_DEC_WB_RegBank_31_3_port, 
      pipeline_RegFile_DEC_WB_RegBank_31_4_port, 
      pipeline_RegFile_DEC_WB_RegBank_31_5_port, 
      pipeline_RegFile_DEC_WB_RegBank_31_6_port, 
      pipeline_RegFile_DEC_WB_RegBank_31_7_port, 
      pipeline_RegFile_DEC_WB_RegBank_31_8_port, 
      pipeline_RegFile_DEC_WB_RegBank_31_9_port, 
      pipeline_RegFile_DEC_WB_RegBank_31_10_port, 
      pipeline_RegFile_DEC_WB_RegBank_31_11_port, 
      pipeline_RegFile_DEC_WB_RegBank_31_12_port, 
      pipeline_RegFile_DEC_WB_RegBank_31_13_port, 
      pipeline_RegFile_DEC_WB_RegBank_31_14_port, 
      pipeline_RegFile_DEC_WB_RegBank_31_15_port, 
      pipeline_RegFile_DEC_WB_RegBank_31_16_port, 
      pipeline_RegFile_DEC_WB_RegBank_31_17_port, 
      pipeline_RegFile_DEC_WB_RegBank_31_18_port, 
      pipeline_RegFile_DEC_WB_RegBank_31_19_port, 
      pipeline_RegFile_DEC_WB_RegBank_31_20_port, 
      pipeline_RegFile_DEC_WB_RegBank_31_21_port, 
      pipeline_RegFile_DEC_WB_RegBank_31_22_port, 
      pipeline_RegFile_DEC_WB_RegBank_31_23_port, 
      pipeline_RegFile_DEC_WB_RegBank_31_24_port, 
      pipeline_RegFile_DEC_WB_RegBank_31_25_port, 
      pipeline_RegFile_DEC_WB_RegBank_31_26_port, 
      pipeline_RegFile_DEC_WB_RegBank_31_27_port, 
      pipeline_RegFile_DEC_WB_RegBank_31_28_port, 
      pipeline_RegFile_DEC_WB_RegBank_31_29_port, 
      pipeline_RegFile_DEC_WB_RegBank_31_30_port, 
      pipeline_RegFile_DEC_WB_RegBank_31_31_port, 
      pipeline_RegFile_DEC_WB_RegBank_30_0_port, 
      pipeline_RegFile_DEC_WB_RegBank_30_1_port, 
      pipeline_RegFile_DEC_WB_RegBank_30_2_port, 
      pipeline_RegFile_DEC_WB_RegBank_30_3_port, 
      pipeline_RegFile_DEC_WB_RegBank_30_4_port, 
      pipeline_RegFile_DEC_WB_RegBank_30_5_port, 
      pipeline_RegFile_DEC_WB_RegBank_30_6_port, 
      pipeline_RegFile_DEC_WB_RegBank_30_7_port, 
      pipeline_RegFile_DEC_WB_RegBank_30_8_port, 
      pipeline_RegFile_DEC_WB_RegBank_30_9_port, 
      pipeline_RegFile_DEC_WB_RegBank_30_10_port, 
      pipeline_RegFile_DEC_WB_RegBank_30_11_port, 
      pipeline_RegFile_DEC_WB_RegBank_30_12_port, 
      pipeline_RegFile_DEC_WB_RegBank_30_13_port, 
      pipeline_RegFile_DEC_WB_RegBank_30_14_port, 
      pipeline_RegFile_DEC_WB_RegBank_30_15_port, 
      pipeline_RegFile_DEC_WB_RegBank_30_16_port, 
      pipeline_RegFile_DEC_WB_RegBank_30_17_port, 
      pipeline_RegFile_DEC_WB_RegBank_30_18_port, 
      pipeline_RegFile_DEC_WB_RegBank_30_19_port, 
      pipeline_RegFile_DEC_WB_RegBank_30_20_port, 
      pipeline_RegFile_DEC_WB_RegBank_30_21_port, 
      pipeline_RegFile_DEC_WB_RegBank_30_22_port, 
      pipeline_RegFile_DEC_WB_RegBank_30_23_port, 
      pipeline_RegFile_DEC_WB_RegBank_30_24_port, 
      pipeline_RegFile_DEC_WB_RegBank_30_25_port, 
      pipeline_RegFile_DEC_WB_RegBank_30_26_port, 
      pipeline_RegFile_DEC_WB_RegBank_30_27_port, 
      pipeline_RegFile_DEC_WB_RegBank_30_28_port, 
      pipeline_RegFile_DEC_WB_RegBank_30_29_port, 
      pipeline_RegFile_DEC_WB_RegBank_30_30_port, 
      pipeline_RegFile_DEC_WB_RegBank_30_31_port, 
      pipeline_RegFile_DEC_WB_RegBank_29_0_port, 
      pipeline_RegFile_DEC_WB_RegBank_29_1_port, 
      pipeline_RegFile_DEC_WB_RegBank_29_2_port, 
      pipeline_RegFile_DEC_WB_RegBank_29_3_port, 
      pipeline_RegFile_DEC_WB_RegBank_29_4_port, 
      pipeline_RegFile_DEC_WB_RegBank_29_5_port, 
      pipeline_RegFile_DEC_WB_RegBank_29_6_port, 
      pipeline_RegFile_DEC_WB_RegBank_29_7_port, 
      pipeline_RegFile_DEC_WB_RegBank_29_8_port, 
      pipeline_RegFile_DEC_WB_RegBank_29_9_port, 
      pipeline_RegFile_DEC_WB_RegBank_29_10_port, 
      pipeline_RegFile_DEC_WB_RegBank_29_11_port, 
      pipeline_RegFile_DEC_WB_RegBank_29_12_port, 
      pipeline_RegFile_DEC_WB_RegBank_29_13_port, 
      pipeline_RegFile_DEC_WB_RegBank_29_14_port, 
      pipeline_RegFile_DEC_WB_RegBank_29_15_port, 
      pipeline_RegFile_DEC_WB_RegBank_29_16_port, 
      pipeline_RegFile_DEC_WB_RegBank_29_17_port, 
      pipeline_RegFile_DEC_WB_RegBank_29_18_port, 
      pipeline_RegFile_DEC_WB_RegBank_29_19_port, 
      pipeline_RegFile_DEC_WB_RegBank_29_20_port, 
      pipeline_RegFile_DEC_WB_RegBank_29_21_port, 
      pipeline_RegFile_DEC_WB_RegBank_29_22_port, 
      pipeline_RegFile_DEC_WB_RegBank_29_23_port, 
      pipeline_RegFile_DEC_WB_RegBank_29_24_port, 
      pipeline_RegFile_DEC_WB_RegBank_29_25_port, 
      pipeline_RegFile_DEC_WB_RegBank_29_26_port, 
      pipeline_RegFile_DEC_WB_RegBank_29_27_port, 
      pipeline_RegFile_DEC_WB_RegBank_29_28_port, 
      pipeline_RegFile_DEC_WB_RegBank_29_29_port, 
      pipeline_RegFile_DEC_WB_RegBank_29_30_port, 
      pipeline_RegFile_DEC_WB_RegBank_29_31_port, 
      pipeline_RegFile_DEC_WB_RegBank_28_0_port, 
      pipeline_RegFile_DEC_WB_RegBank_28_1_port, 
      pipeline_RegFile_DEC_WB_RegBank_28_2_port, 
      pipeline_RegFile_DEC_WB_RegBank_28_3_port, 
      pipeline_RegFile_DEC_WB_RegBank_28_4_port, 
      pipeline_RegFile_DEC_WB_RegBank_28_5_port, 
      pipeline_RegFile_DEC_WB_RegBank_28_6_port, 
      pipeline_RegFile_DEC_WB_RegBank_28_7_port, 
      pipeline_RegFile_DEC_WB_RegBank_28_8_port, 
      pipeline_RegFile_DEC_WB_RegBank_28_9_port, 
      pipeline_RegFile_DEC_WB_RegBank_28_10_port, 
      pipeline_RegFile_DEC_WB_RegBank_28_11_port, 
      pipeline_RegFile_DEC_WB_RegBank_28_12_port, 
      pipeline_RegFile_DEC_WB_RegBank_28_13_port, 
      pipeline_RegFile_DEC_WB_RegBank_28_14_port, 
      pipeline_RegFile_DEC_WB_RegBank_28_15_port, 
      pipeline_RegFile_DEC_WB_RegBank_28_16_port, 
      pipeline_RegFile_DEC_WB_RegBank_28_17_port, 
      pipeline_RegFile_DEC_WB_RegBank_28_18_port, 
      pipeline_RegFile_DEC_WB_RegBank_28_19_port, 
      pipeline_RegFile_DEC_WB_RegBank_28_20_port, 
      pipeline_RegFile_DEC_WB_RegBank_28_21_port, 
      pipeline_RegFile_DEC_WB_RegBank_28_22_port, 
      pipeline_RegFile_DEC_WB_RegBank_28_23_port, 
      pipeline_RegFile_DEC_WB_RegBank_28_24_port, 
      pipeline_RegFile_DEC_WB_RegBank_28_25_port, 
      pipeline_RegFile_DEC_WB_RegBank_28_26_port, 
      pipeline_RegFile_DEC_WB_RegBank_28_27_port, 
      pipeline_RegFile_DEC_WB_RegBank_28_28_port, 
      pipeline_RegFile_DEC_WB_RegBank_28_29_port, 
      pipeline_RegFile_DEC_WB_RegBank_28_30_port, 
      pipeline_RegFile_DEC_WB_RegBank_28_31_port, 
      pipeline_RegFile_DEC_WB_RegBank_27_0_port, 
      pipeline_RegFile_DEC_WB_RegBank_27_1_port, 
      pipeline_RegFile_DEC_WB_RegBank_27_2_port, 
      pipeline_RegFile_DEC_WB_RegBank_27_3_port, 
      pipeline_RegFile_DEC_WB_RegBank_27_4_port, 
      pipeline_RegFile_DEC_WB_RegBank_27_5_port, 
      pipeline_RegFile_DEC_WB_RegBank_27_6_port, 
      pipeline_RegFile_DEC_WB_RegBank_27_7_port, 
      pipeline_RegFile_DEC_WB_RegBank_27_8_port, 
      pipeline_RegFile_DEC_WB_RegBank_27_9_port, 
      pipeline_RegFile_DEC_WB_RegBank_27_10_port, 
      pipeline_RegFile_DEC_WB_RegBank_27_11_port, 
      pipeline_RegFile_DEC_WB_RegBank_27_12_port, 
      pipeline_RegFile_DEC_WB_RegBank_27_13_port, 
      pipeline_RegFile_DEC_WB_RegBank_27_14_port, 
      pipeline_RegFile_DEC_WB_RegBank_27_15_port, 
      pipeline_RegFile_DEC_WB_RegBank_27_16_port, 
      pipeline_RegFile_DEC_WB_RegBank_27_17_port, 
      pipeline_RegFile_DEC_WB_RegBank_27_18_port, 
      pipeline_RegFile_DEC_WB_RegBank_27_19_port, 
      pipeline_RegFile_DEC_WB_RegBank_27_20_port, 
      pipeline_RegFile_DEC_WB_RegBank_27_21_port, 
      pipeline_RegFile_DEC_WB_RegBank_27_22_port, 
      pipeline_RegFile_DEC_WB_RegBank_27_23_port, 
      pipeline_RegFile_DEC_WB_RegBank_27_24_port, 
      pipeline_RegFile_DEC_WB_RegBank_27_25_port, 
      pipeline_RegFile_DEC_WB_RegBank_27_26_port, 
      pipeline_RegFile_DEC_WB_RegBank_27_27_port, 
      pipeline_RegFile_DEC_WB_RegBank_27_28_port, 
      pipeline_RegFile_DEC_WB_RegBank_27_29_port, 
      pipeline_RegFile_DEC_WB_RegBank_27_30_port, 
      pipeline_RegFile_DEC_WB_RegBank_27_31_port, 
      pipeline_RegFile_DEC_WB_RegBank_26_0_port, 
      pipeline_RegFile_DEC_WB_RegBank_26_1_port, 
      pipeline_RegFile_DEC_WB_RegBank_26_2_port, 
      pipeline_RegFile_DEC_WB_RegBank_26_3_port, 
      pipeline_RegFile_DEC_WB_RegBank_26_4_port, 
      pipeline_RegFile_DEC_WB_RegBank_26_5_port, 
      pipeline_RegFile_DEC_WB_RegBank_26_6_port, 
      pipeline_RegFile_DEC_WB_RegBank_26_7_port, 
      pipeline_RegFile_DEC_WB_RegBank_26_8_port, 
      pipeline_RegFile_DEC_WB_RegBank_26_9_port, 
      pipeline_RegFile_DEC_WB_RegBank_26_10_port, 
      pipeline_RegFile_DEC_WB_RegBank_26_11_port, 
      pipeline_RegFile_DEC_WB_RegBank_26_12_port, 
      pipeline_RegFile_DEC_WB_RegBank_26_13_port, 
      pipeline_RegFile_DEC_WB_RegBank_26_14_port, 
      pipeline_RegFile_DEC_WB_RegBank_26_15_port, 
      pipeline_RegFile_DEC_WB_RegBank_26_16_port, 
      pipeline_RegFile_DEC_WB_RegBank_26_17_port, 
      pipeline_RegFile_DEC_WB_RegBank_26_18_port, 
      pipeline_RegFile_DEC_WB_RegBank_26_19_port, 
      pipeline_RegFile_DEC_WB_RegBank_26_20_port, 
      pipeline_RegFile_DEC_WB_RegBank_26_21_port, 
      pipeline_RegFile_DEC_WB_RegBank_26_22_port, 
      pipeline_RegFile_DEC_WB_RegBank_26_23_port, 
      pipeline_RegFile_DEC_WB_RegBank_26_24_port, 
      pipeline_RegFile_DEC_WB_RegBank_26_25_port, 
      pipeline_RegFile_DEC_WB_RegBank_26_26_port, 
      pipeline_RegFile_DEC_WB_RegBank_26_27_port, 
      pipeline_RegFile_DEC_WB_RegBank_26_28_port, 
      pipeline_RegFile_DEC_WB_RegBank_26_29_port, 
      pipeline_RegFile_DEC_WB_RegBank_26_30_port, 
      pipeline_RegFile_DEC_WB_RegBank_26_31_port, 
      pipeline_RegFile_DEC_WB_RegBank_25_0_port, 
      pipeline_RegFile_DEC_WB_RegBank_25_1_port, 
      pipeline_RegFile_DEC_WB_RegBank_25_2_port, 
      pipeline_RegFile_DEC_WB_RegBank_25_3_port, 
      pipeline_RegFile_DEC_WB_RegBank_25_4_port, 
      pipeline_RegFile_DEC_WB_RegBank_25_5_port, 
      pipeline_RegFile_DEC_WB_RegBank_25_6_port, 
      pipeline_RegFile_DEC_WB_RegBank_25_7_port, 
      pipeline_RegFile_DEC_WB_RegBank_25_8_port, 
      pipeline_RegFile_DEC_WB_RegBank_25_9_port, 
      pipeline_RegFile_DEC_WB_RegBank_25_10_port, 
      pipeline_RegFile_DEC_WB_RegBank_25_11_port, 
      pipeline_RegFile_DEC_WB_RegBank_25_12_port, 
      pipeline_RegFile_DEC_WB_RegBank_25_13_port, 
      pipeline_RegFile_DEC_WB_RegBank_25_14_port, 
      pipeline_RegFile_DEC_WB_RegBank_25_15_port, 
      pipeline_RegFile_DEC_WB_RegBank_25_16_port, 
      pipeline_RegFile_DEC_WB_RegBank_25_17_port, 
      pipeline_RegFile_DEC_WB_RegBank_25_18_port, 
      pipeline_RegFile_DEC_WB_RegBank_25_19_port, 
      pipeline_RegFile_DEC_WB_RegBank_25_20_port, 
      pipeline_RegFile_DEC_WB_RegBank_25_21_port, 
      pipeline_RegFile_DEC_WB_RegBank_25_22_port, 
      pipeline_RegFile_DEC_WB_RegBank_25_23_port, 
      pipeline_RegFile_DEC_WB_RegBank_25_24_port, 
      pipeline_RegFile_DEC_WB_RegBank_25_25_port, 
      pipeline_RegFile_DEC_WB_RegBank_25_26_port, 
      pipeline_RegFile_DEC_WB_RegBank_25_27_port, 
      pipeline_RegFile_DEC_WB_RegBank_25_28_port, 
      pipeline_RegFile_DEC_WB_RegBank_25_29_port, 
      pipeline_RegFile_DEC_WB_RegBank_25_30_port, 
      pipeline_RegFile_DEC_WB_RegBank_25_31_port, 
      pipeline_RegFile_DEC_WB_RegBank_24_0_port, 
      pipeline_RegFile_DEC_WB_RegBank_24_1_port, 
      pipeline_RegFile_DEC_WB_RegBank_24_2_port, 
      pipeline_RegFile_DEC_WB_RegBank_24_3_port, 
      pipeline_RegFile_DEC_WB_RegBank_24_4_port, 
      pipeline_RegFile_DEC_WB_RegBank_24_5_port, 
      pipeline_RegFile_DEC_WB_RegBank_24_6_port, 
      pipeline_RegFile_DEC_WB_RegBank_24_7_port, 
      pipeline_RegFile_DEC_WB_RegBank_24_8_port, 
      pipeline_RegFile_DEC_WB_RegBank_24_9_port, 
      pipeline_RegFile_DEC_WB_RegBank_24_10_port, 
      pipeline_RegFile_DEC_WB_RegBank_24_11_port, 
      pipeline_RegFile_DEC_WB_RegBank_24_12_port, 
      pipeline_RegFile_DEC_WB_RegBank_24_13_port, 
      pipeline_RegFile_DEC_WB_RegBank_24_14_port, 
      pipeline_RegFile_DEC_WB_RegBank_24_15_port, 
      pipeline_RegFile_DEC_WB_RegBank_24_16_port, 
      pipeline_RegFile_DEC_WB_RegBank_24_17_port, 
      pipeline_RegFile_DEC_WB_RegBank_24_18_port, 
      pipeline_RegFile_DEC_WB_RegBank_24_19_port, 
      pipeline_RegFile_DEC_WB_RegBank_24_20_port, 
      pipeline_RegFile_DEC_WB_RegBank_24_21_port, 
      pipeline_RegFile_DEC_WB_RegBank_24_22_port, 
      pipeline_RegFile_DEC_WB_RegBank_24_23_port, 
      pipeline_RegFile_DEC_WB_RegBank_24_24_port, 
      pipeline_RegFile_DEC_WB_RegBank_24_25_port, 
      pipeline_RegFile_DEC_WB_RegBank_24_26_port, 
      pipeline_RegFile_DEC_WB_RegBank_24_27_port, 
      pipeline_RegFile_DEC_WB_RegBank_24_28_port, 
      pipeline_RegFile_DEC_WB_RegBank_24_29_port, 
      pipeline_RegFile_DEC_WB_RegBank_24_30_port, 
      pipeline_RegFile_DEC_WB_RegBank_24_31_port, 
      pipeline_RegFile_DEC_WB_RegBank_23_0_port, 
      pipeline_RegFile_DEC_WB_RegBank_23_1_port, 
      pipeline_RegFile_DEC_WB_RegBank_23_2_port, 
      pipeline_RegFile_DEC_WB_RegBank_23_3_port, 
      pipeline_RegFile_DEC_WB_RegBank_23_4_port, 
      pipeline_RegFile_DEC_WB_RegBank_23_5_port, 
      pipeline_RegFile_DEC_WB_RegBank_23_6_port, 
      pipeline_RegFile_DEC_WB_RegBank_23_7_port, 
      pipeline_RegFile_DEC_WB_RegBank_23_8_port, 
      pipeline_RegFile_DEC_WB_RegBank_23_9_port, 
      pipeline_RegFile_DEC_WB_RegBank_23_10_port, 
      pipeline_RegFile_DEC_WB_RegBank_23_11_port, 
      pipeline_RegFile_DEC_WB_RegBank_23_12_port, 
      pipeline_RegFile_DEC_WB_RegBank_23_13_port, 
      pipeline_RegFile_DEC_WB_RegBank_23_14_port, 
      pipeline_RegFile_DEC_WB_RegBank_23_15_port, 
      pipeline_RegFile_DEC_WB_RegBank_23_16_port, 
      pipeline_RegFile_DEC_WB_RegBank_23_17_port, 
      pipeline_RegFile_DEC_WB_RegBank_23_18_port, 
      pipeline_RegFile_DEC_WB_RegBank_23_19_port, 
      pipeline_RegFile_DEC_WB_RegBank_23_20_port, 
      pipeline_RegFile_DEC_WB_RegBank_23_21_port, 
      pipeline_RegFile_DEC_WB_RegBank_23_22_port, 
      pipeline_RegFile_DEC_WB_RegBank_23_23_port, 
      pipeline_RegFile_DEC_WB_RegBank_23_24_port, 
      pipeline_RegFile_DEC_WB_RegBank_23_25_port, 
      pipeline_RegFile_DEC_WB_RegBank_23_26_port, 
      pipeline_RegFile_DEC_WB_RegBank_23_27_port, 
      pipeline_RegFile_DEC_WB_RegBank_23_28_port, 
      pipeline_RegFile_DEC_WB_RegBank_23_29_port, 
      pipeline_RegFile_DEC_WB_RegBank_23_30_port, 
      pipeline_RegFile_DEC_WB_RegBank_23_31_port, 
      pipeline_RegFile_DEC_WB_RegBank_22_0_port, 
      pipeline_RegFile_DEC_WB_RegBank_22_1_port, 
      pipeline_RegFile_DEC_WB_RegBank_22_2_port, 
      pipeline_RegFile_DEC_WB_RegBank_22_3_port, 
      pipeline_RegFile_DEC_WB_RegBank_22_4_port, 
      pipeline_RegFile_DEC_WB_RegBank_22_5_port, 
      pipeline_RegFile_DEC_WB_RegBank_22_6_port, 
      pipeline_RegFile_DEC_WB_RegBank_22_7_port, 
      pipeline_RegFile_DEC_WB_RegBank_22_8_port, 
      pipeline_RegFile_DEC_WB_RegBank_22_9_port, 
      pipeline_RegFile_DEC_WB_RegBank_22_10_port, 
      pipeline_RegFile_DEC_WB_RegBank_22_11_port, 
      pipeline_RegFile_DEC_WB_RegBank_22_12_port, 
      pipeline_RegFile_DEC_WB_RegBank_22_13_port, 
      pipeline_RegFile_DEC_WB_RegBank_22_14_port, 
      pipeline_RegFile_DEC_WB_RegBank_22_15_port, 
      pipeline_RegFile_DEC_WB_RegBank_22_16_port, 
      pipeline_RegFile_DEC_WB_RegBank_22_17_port, 
      pipeline_RegFile_DEC_WB_RegBank_22_18_port, 
      pipeline_RegFile_DEC_WB_RegBank_22_19_port, 
      pipeline_RegFile_DEC_WB_RegBank_22_20_port, 
      pipeline_RegFile_DEC_WB_RegBank_22_21_port, 
      pipeline_RegFile_DEC_WB_RegBank_22_22_port, 
      pipeline_RegFile_DEC_WB_RegBank_22_23_port, 
      pipeline_RegFile_DEC_WB_RegBank_22_24_port, 
      pipeline_RegFile_DEC_WB_RegBank_22_25_port, 
      pipeline_RegFile_DEC_WB_RegBank_22_26_port, 
      pipeline_RegFile_DEC_WB_RegBank_22_27_port, 
      pipeline_RegFile_DEC_WB_RegBank_22_28_port, 
      pipeline_RegFile_DEC_WB_RegBank_22_29_port, 
      pipeline_RegFile_DEC_WB_RegBank_22_30_port, 
      pipeline_RegFile_DEC_WB_RegBank_22_31_port, 
      pipeline_RegFile_DEC_WB_RegBank_21_0_port, 
      pipeline_RegFile_DEC_WB_RegBank_21_1_port, 
      pipeline_RegFile_DEC_WB_RegBank_21_2_port, 
      pipeline_RegFile_DEC_WB_RegBank_21_3_port, 
      pipeline_RegFile_DEC_WB_RegBank_21_4_port, 
      pipeline_RegFile_DEC_WB_RegBank_21_5_port, 
      pipeline_RegFile_DEC_WB_RegBank_21_6_port, 
      pipeline_RegFile_DEC_WB_RegBank_21_7_port, 
      pipeline_RegFile_DEC_WB_RegBank_21_8_port, 
      pipeline_RegFile_DEC_WB_RegBank_21_9_port, 
      pipeline_RegFile_DEC_WB_RegBank_21_10_port, 
      pipeline_RegFile_DEC_WB_RegBank_21_11_port, 
      pipeline_RegFile_DEC_WB_RegBank_21_12_port, 
      pipeline_RegFile_DEC_WB_RegBank_21_13_port, 
      pipeline_RegFile_DEC_WB_RegBank_21_14_port, 
      pipeline_RegFile_DEC_WB_RegBank_21_15_port, 
      pipeline_RegFile_DEC_WB_RegBank_21_16_port, 
      pipeline_RegFile_DEC_WB_RegBank_21_17_port, 
      pipeline_RegFile_DEC_WB_RegBank_21_18_port, 
      pipeline_RegFile_DEC_WB_RegBank_21_19_port, 
      pipeline_RegFile_DEC_WB_RegBank_21_20_port, 
      pipeline_RegFile_DEC_WB_RegBank_21_21_port, 
      pipeline_RegFile_DEC_WB_RegBank_21_22_port, 
      pipeline_RegFile_DEC_WB_RegBank_21_23_port, 
      pipeline_RegFile_DEC_WB_RegBank_21_24_port, 
      pipeline_RegFile_DEC_WB_RegBank_21_25_port, 
      pipeline_RegFile_DEC_WB_RegBank_21_26_port, 
      pipeline_RegFile_DEC_WB_RegBank_21_27_port, 
      pipeline_RegFile_DEC_WB_RegBank_21_28_port, 
      pipeline_RegFile_DEC_WB_RegBank_21_29_port, 
      pipeline_RegFile_DEC_WB_RegBank_21_30_port, 
      pipeline_RegFile_DEC_WB_RegBank_21_31_port, 
      pipeline_RegFile_DEC_WB_RegBank_20_0_port, 
      pipeline_RegFile_DEC_WB_RegBank_20_1_port, 
      pipeline_RegFile_DEC_WB_RegBank_20_2_port, 
      pipeline_RegFile_DEC_WB_RegBank_20_3_port, 
      pipeline_RegFile_DEC_WB_RegBank_20_4_port, 
      pipeline_RegFile_DEC_WB_RegBank_20_5_port, 
      pipeline_RegFile_DEC_WB_RegBank_20_6_port, 
      pipeline_RegFile_DEC_WB_RegBank_20_7_port, 
      pipeline_RegFile_DEC_WB_RegBank_20_8_port, 
      pipeline_RegFile_DEC_WB_RegBank_20_9_port, 
      pipeline_RegFile_DEC_WB_RegBank_20_10_port, 
      pipeline_RegFile_DEC_WB_RegBank_20_11_port, 
      pipeline_RegFile_DEC_WB_RegBank_20_12_port, 
      pipeline_RegFile_DEC_WB_RegBank_20_13_port, 
      pipeline_RegFile_DEC_WB_RegBank_20_14_port, 
      pipeline_RegFile_DEC_WB_RegBank_20_15_port, 
      pipeline_RegFile_DEC_WB_RegBank_20_16_port, 
      pipeline_RegFile_DEC_WB_RegBank_20_17_port, 
      pipeline_RegFile_DEC_WB_RegBank_20_18_port, 
      pipeline_RegFile_DEC_WB_RegBank_20_19_port, 
      pipeline_RegFile_DEC_WB_RegBank_20_20_port, 
      pipeline_RegFile_DEC_WB_RegBank_20_21_port, 
      pipeline_RegFile_DEC_WB_RegBank_20_22_port, 
      pipeline_RegFile_DEC_WB_RegBank_20_23_port, 
      pipeline_RegFile_DEC_WB_RegBank_20_24_port, 
      pipeline_RegFile_DEC_WB_RegBank_20_25_port, 
      pipeline_RegFile_DEC_WB_RegBank_20_26_port, 
      pipeline_RegFile_DEC_WB_RegBank_20_27_port, 
      pipeline_RegFile_DEC_WB_RegBank_20_28_port, 
      pipeline_RegFile_DEC_WB_RegBank_20_29_port, 
      pipeline_RegFile_DEC_WB_RegBank_20_30_port, 
      pipeline_RegFile_DEC_WB_RegBank_20_31_port, 
      pipeline_RegFile_DEC_WB_RegBank_19_0_port, 
      pipeline_RegFile_DEC_WB_RegBank_19_1_port, 
      pipeline_RegFile_DEC_WB_RegBank_19_2_port, 
      pipeline_RegFile_DEC_WB_RegBank_19_3_port, 
      pipeline_RegFile_DEC_WB_RegBank_19_4_port, 
      pipeline_RegFile_DEC_WB_RegBank_19_5_port, 
      pipeline_RegFile_DEC_WB_RegBank_19_6_port, 
      pipeline_RegFile_DEC_WB_RegBank_19_7_port, 
      pipeline_RegFile_DEC_WB_RegBank_19_8_port, 
      pipeline_RegFile_DEC_WB_RegBank_19_9_port, 
      pipeline_RegFile_DEC_WB_RegBank_19_10_port, 
      pipeline_RegFile_DEC_WB_RegBank_19_11_port, 
      pipeline_RegFile_DEC_WB_RegBank_19_12_port, 
      pipeline_RegFile_DEC_WB_RegBank_19_13_port, 
      pipeline_RegFile_DEC_WB_RegBank_19_14_port, 
      pipeline_RegFile_DEC_WB_RegBank_19_15_port, 
      pipeline_RegFile_DEC_WB_RegBank_19_16_port, 
      pipeline_RegFile_DEC_WB_RegBank_19_17_port, 
      pipeline_RegFile_DEC_WB_RegBank_19_18_port, 
      pipeline_RegFile_DEC_WB_RegBank_19_19_port, 
      pipeline_RegFile_DEC_WB_RegBank_19_20_port, 
      pipeline_RegFile_DEC_WB_RegBank_19_21_port, 
      pipeline_RegFile_DEC_WB_RegBank_19_22_port, 
      pipeline_RegFile_DEC_WB_RegBank_19_23_port, 
      pipeline_RegFile_DEC_WB_RegBank_19_24_port, 
      pipeline_RegFile_DEC_WB_RegBank_19_25_port, 
      pipeline_RegFile_DEC_WB_RegBank_19_26_port, 
      pipeline_RegFile_DEC_WB_RegBank_19_27_port, 
      pipeline_RegFile_DEC_WB_RegBank_19_28_port, 
      pipeline_RegFile_DEC_WB_RegBank_19_29_port, 
      pipeline_RegFile_DEC_WB_RegBank_19_30_port, 
      pipeline_RegFile_DEC_WB_RegBank_19_31_port, 
      pipeline_RegFile_DEC_WB_RegBank_18_0_port, 
      pipeline_RegFile_DEC_WB_RegBank_18_1_port, 
      pipeline_RegFile_DEC_WB_RegBank_18_2_port, 
      pipeline_RegFile_DEC_WB_RegBank_18_3_port, 
      pipeline_RegFile_DEC_WB_RegBank_18_4_port, 
      pipeline_RegFile_DEC_WB_RegBank_18_5_port, 
      pipeline_RegFile_DEC_WB_RegBank_18_6_port, 
      pipeline_RegFile_DEC_WB_RegBank_18_7_port, 
      pipeline_RegFile_DEC_WB_RegBank_18_8_port, 
      pipeline_RegFile_DEC_WB_RegBank_18_9_port, 
      pipeline_RegFile_DEC_WB_RegBank_18_10_port, 
      pipeline_RegFile_DEC_WB_RegBank_18_11_port, 
      pipeline_RegFile_DEC_WB_RegBank_18_12_port, 
      pipeline_RegFile_DEC_WB_RegBank_18_13_port, 
      pipeline_RegFile_DEC_WB_RegBank_18_14_port, 
      pipeline_RegFile_DEC_WB_RegBank_18_15_port, 
      pipeline_RegFile_DEC_WB_RegBank_18_16_port, 
      pipeline_RegFile_DEC_WB_RegBank_18_17_port, 
      pipeline_RegFile_DEC_WB_RegBank_18_18_port, 
      pipeline_RegFile_DEC_WB_RegBank_18_19_port, 
      pipeline_RegFile_DEC_WB_RegBank_18_20_port, 
      pipeline_RegFile_DEC_WB_RegBank_18_21_port, 
      pipeline_RegFile_DEC_WB_RegBank_18_22_port, 
      pipeline_RegFile_DEC_WB_RegBank_18_23_port, 
      pipeline_RegFile_DEC_WB_RegBank_18_24_port, 
      pipeline_RegFile_DEC_WB_RegBank_18_25_port, 
      pipeline_RegFile_DEC_WB_RegBank_18_26_port, 
      pipeline_RegFile_DEC_WB_RegBank_18_27_port, 
      pipeline_RegFile_DEC_WB_RegBank_18_28_port, 
      pipeline_RegFile_DEC_WB_RegBank_18_29_port, 
      pipeline_RegFile_DEC_WB_RegBank_18_30_port, 
      pipeline_RegFile_DEC_WB_RegBank_18_31_port, 
      pipeline_RegFile_DEC_WB_RegBank_17_0_port, 
      pipeline_RegFile_DEC_WB_RegBank_17_1_port, 
      pipeline_RegFile_DEC_WB_RegBank_17_2_port, 
      pipeline_RegFile_DEC_WB_RegBank_17_3_port, 
      pipeline_RegFile_DEC_WB_RegBank_17_4_port, 
      pipeline_RegFile_DEC_WB_RegBank_17_5_port, 
      pipeline_RegFile_DEC_WB_RegBank_17_6_port, 
      pipeline_RegFile_DEC_WB_RegBank_17_7_port, 
      pipeline_RegFile_DEC_WB_RegBank_17_8_port, 
      pipeline_RegFile_DEC_WB_RegBank_17_9_port, 
      pipeline_RegFile_DEC_WB_RegBank_17_10_port, 
      pipeline_RegFile_DEC_WB_RegBank_17_11_port, 
      pipeline_RegFile_DEC_WB_RegBank_17_12_port, 
      pipeline_RegFile_DEC_WB_RegBank_17_13_port, 
      pipeline_RegFile_DEC_WB_RegBank_17_14_port, 
      pipeline_RegFile_DEC_WB_RegBank_17_15_port, 
      pipeline_RegFile_DEC_WB_RegBank_17_16_port, 
      pipeline_RegFile_DEC_WB_RegBank_17_17_port, 
      pipeline_RegFile_DEC_WB_RegBank_17_18_port, 
      pipeline_RegFile_DEC_WB_RegBank_17_19_port, 
      pipeline_RegFile_DEC_WB_RegBank_17_20_port, 
      pipeline_RegFile_DEC_WB_RegBank_17_21_port, 
      pipeline_RegFile_DEC_WB_RegBank_17_22_port, 
      pipeline_RegFile_DEC_WB_RegBank_17_23_port, 
      pipeline_RegFile_DEC_WB_RegBank_17_24_port, 
      pipeline_RegFile_DEC_WB_RegBank_17_25_port, 
      pipeline_RegFile_DEC_WB_RegBank_17_26_port, 
      pipeline_RegFile_DEC_WB_RegBank_17_27_port, 
      pipeline_RegFile_DEC_WB_RegBank_17_28_port, 
      pipeline_RegFile_DEC_WB_RegBank_17_29_port, 
      pipeline_RegFile_DEC_WB_RegBank_17_30_port, 
      pipeline_RegFile_DEC_WB_RegBank_17_31_port, 
      pipeline_RegFile_DEC_WB_RegBank_16_0_port, 
      pipeline_RegFile_DEC_WB_RegBank_16_1_port, 
      pipeline_RegFile_DEC_WB_RegBank_16_2_port, 
      pipeline_RegFile_DEC_WB_RegBank_16_3_port, 
      pipeline_RegFile_DEC_WB_RegBank_16_4_port, 
      pipeline_RegFile_DEC_WB_RegBank_16_5_port, 
      pipeline_RegFile_DEC_WB_RegBank_16_6_port, 
      pipeline_RegFile_DEC_WB_RegBank_16_7_port, 
      pipeline_RegFile_DEC_WB_RegBank_16_8_port, 
      pipeline_RegFile_DEC_WB_RegBank_16_9_port, 
      pipeline_RegFile_DEC_WB_RegBank_16_10_port, 
      pipeline_RegFile_DEC_WB_RegBank_16_11_port, 
      pipeline_RegFile_DEC_WB_RegBank_16_12_port, 
      pipeline_RegFile_DEC_WB_RegBank_16_13_port, 
      pipeline_RegFile_DEC_WB_RegBank_16_14_port, 
      pipeline_RegFile_DEC_WB_RegBank_16_15_port, 
      pipeline_RegFile_DEC_WB_RegBank_16_16_port, 
      pipeline_RegFile_DEC_WB_RegBank_16_17_port, 
      pipeline_RegFile_DEC_WB_RegBank_16_18_port, 
      pipeline_RegFile_DEC_WB_RegBank_16_19_port, 
      pipeline_RegFile_DEC_WB_RegBank_16_20_port, 
      pipeline_RegFile_DEC_WB_RegBank_16_21_port, 
      pipeline_RegFile_DEC_WB_RegBank_16_22_port, 
      pipeline_RegFile_DEC_WB_RegBank_16_23_port, 
      pipeline_RegFile_DEC_WB_RegBank_16_24_port, 
      pipeline_RegFile_DEC_WB_RegBank_16_25_port, 
      pipeline_RegFile_DEC_WB_RegBank_16_26_port, 
      pipeline_RegFile_DEC_WB_RegBank_16_27_port, 
      pipeline_RegFile_DEC_WB_RegBank_16_28_port, 
      pipeline_RegFile_DEC_WB_RegBank_16_29_port, 
      pipeline_RegFile_DEC_WB_RegBank_16_30_port, 
      pipeline_RegFile_DEC_WB_RegBank_16_31_port, 
      pipeline_RegFile_DEC_WB_RegBank_15_0_port, 
      pipeline_RegFile_DEC_WB_RegBank_15_1_port, 
      pipeline_RegFile_DEC_WB_RegBank_15_2_port, 
      pipeline_RegFile_DEC_WB_RegBank_15_3_port, 
      pipeline_RegFile_DEC_WB_RegBank_15_4_port, 
      pipeline_RegFile_DEC_WB_RegBank_15_5_port, 
      pipeline_RegFile_DEC_WB_RegBank_15_6_port, 
      pipeline_RegFile_DEC_WB_RegBank_15_7_port, 
      pipeline_RegFile_DEC_WB_RegBank_15_8_port, 
      pipeline_RegFile_DEC_WB_RegBank_15_9_port, 
      pipeline_RegFile_DEC_WB_RegBank_15_10_port, 
      pipeline_RegFile_DEC_WB_RegBank_15_11_port, 
      pipeline_RegFile_DEC_WB_RegBank_15_12_port, 
      pipeline_RegFile_DEC_WB_RegBank_15_13_port, 
      pipeline_RegFile_DEC_WB_RegBank_15_14_port, 
      pipeline_RegFile_DEC_WB_RegBank_15_15_port, 
      pipeline_RegFile_DEC_WB_RegBank_15_16_port, 
      pipeline_RegFile_DEC_WB_RegBank_15_17_port, 
      pipeline_RegFile_DEC_WB_RegBank_15_18_port, 
      pipeline_RegFile_DEC_WB_RegBank_15_19_port, 
      pipeline_RegFile_DEC_WB_RegBank_15_20_port, 
      pipeline_RegFile_DEC_WB_RegBank_15_21_port, 
      pipeline_RegFile_DEC_WB_RegBank_15_22_port, 
      pipeline_RegFile_DEC_WB_RegBank_15_23_port, 
      pipeline_RegFile_DEC_WB_RegBank_15_24_port, 
      pipeline_RegFile_DEC_WB_RegBank_15_25_port, 
      pipeline_RegFile_DEC_WB_RegBank_15_26_port, 
      pipeline_RegFile_DEC_WB_RegBank_15_27_port, 
      pipeline_RegFile_DEC_WB_RegBank_15_28_port, 
      pipeline_RegFile_DEC_WB_RegBank_15_29_port, 
      pipeline_RegFile_DEC_WB_RegBank_15_30_port, 
      pipeline_RegFile_DEC_WB_RegBank_15_31_port, 
      pipeline_RegFile_DEC_WB_RegBank_14_0_port, 
      pipeline_RegFile_DEC_WB_RegBank_14_1_port, 
      pipeline_RegFile_DEC_WB_RegBank_14_2_port, 
      pipeline_RegFile_DEC_WB_RegBank_14_3_port, 
      pipeline_RegFile_DEC_WB_RegBank_14_4_port, 
      pipeline_RegFile_DEC_WB_RegBank_14_5_port, 
      pipeline_RegFile_DEC_WB_RegBank_14_6_port, 
      pipeline_RegFile_DEC_WB_RegBank_14_7_port, 
      pipeline_RegFile_DEC_WB_RegBank_14_8_port, 
      pipeline_RegFile_DEC_WB_RegBank_14_9_port, 
      pipeline_RegFile_DEC_WB_RegBank_14_10_port, 
      pipeline_RegFile_DEC_WB_RegBank_14_11_port, 
      pipeline_RegFile_DEC_WB_RegBank_14_12_port, 
      pipeline_RegFile_DEC_WB_RegBank_14_13_port, 
      pipeline_RegFile_DEC_WB_RegBank_14_14_port, 
      pipeline_RegFile_DEC_WB_RegBank_14_15_port, 
      pipeline_RegFile_DEC_WB_RegBank_14_16_port, 
      pipeline_RegFile_DEC_WB_RegBank_14_17_port, 
      pipeline_RegFile_DEC_WB_RegBank_14_18_port, 
      pipeline_RegFile_DEC_WB_RegBank_14_19_port, 
      pipeline_RegFile_DEC_WB_RegBank_14_20_port, 
      pipeline_RegFile_DEC_WB_RegBank_14_21_port, 
      pipeline_RegFile_DEC_WB_RegBank_14_22_port, 
      pipeline_RegFile_DEC_WB_RegBank_14_23_port, 
      pipeline_RegFile_DEC_WB_RegBank_14_24_port, 
      pipeline_RegFile_DEC_WB_RegBank_14_25_port, 
      pipeline_RegFile_DEC_WB_RegBank_14_26_port, 
      pipeline_RegFile_DEC_WB_RegBank_14_27_port, 
      pipeline_RegFile_DEC_WB_RegBank_14_28_port, 
      pipeline_RegFile_DEC_WB_RegBank_14_29_port, 
      pipeline_RegFile_DEC_WB_RegBank_14_30_port, 
      pipeline_RegFile_DEC_WB_RegBank_14_31_port, 
      pipeline_RegFile_DEC_WB_RegBank_13_0_port, 
      pipeline_RegFile_DEC_WB_RegBank_13_1_port, 
      pipeline_RegFile_DEC_WB_RegBank_13_2_port, 
      pipeline_RegFile_DEC_WB_RegBank_13_3_port, 
      pipeline_RegFile_DEC_WB_RegBank_13_4_port, 
      pipeline_RegFile_DEC_WB_RegBank_13_5_port, 
      pipeline_RegFile_DEC_WB_RegBank_13_6_port, 
      pipeline_RegFile_DEC_WB_RegBank_13_7_port, 
      pipeline_RegFile_DEC_WB_RegBank_13_8_port, 
      pipeline_RegFile_DEC_WB_RegBank_13_9_port, 
      pipeline_RegFile_DEC_WB_RegBank_13_10_port, 
      pipeline_RegFile_DEC_WB_RegBank_13_11_port, 
      pipeline_RegFile_DEC_WB_RegBank_13_12_port, 
      pipeline_RegFile_DEC_WB_RegBank_13_13_port, 
      pipeline_RegFile_DEC_WB_RegBank_13_14_port, 
      pipeline_RegFile_DEC_WB_RegBank_13_15_port, 
      pipeline_RegFile_DEC_WB_RegBank_13_16_port, 
      pipeline_RegFile_DEC_WB_RegBank_13_17_port, 
      pipeline_RegFile_DEC_WB_RegBank_13_18_port, 
      pipeline_RegFile_DEC_WB_RegBank_13_19_port, 
      pipeline_RegFile_DEC_WB_RegBank_13_20_port, 
      pipeline_RegFile_DEC_WB_RegBank_13_21_port, 
      pipeline_RegFile_DEC_WB_RegBank_13_22_port, 
      pipeline_RegFile_DEC_WB_RegBank_13_23_port, 
      pipeline_RegFile_DEC_WB_RegBank_13_24_port, 
      pipeline_RegFile_DEC_WB_RegBank_13_25_port, 
      pipeline_RegFile_DEC_WB_RegBank_13_26_port, 
      pipeline_RegFile_DEC_WB_RegBank_13_27_port, 
      pipeline_RegFile_DEC_WB_RegBank_13_28_port, 
      pipeline_RegFile_DEC_WB_RegBank_13_29_port, 
      pipeline_RegFile_DEC_WB_RegBank_13_30_port, 
      pipeline_RegFile_DEC_WB_RegBank_13_31_port, 
      pipeline_RegFile_DEC_WB_RegBank_12_0_port, 
      pipeline_RegFile_DEC_WB_RegBank_12_1_port, 
      pipeline_RegFile_DEC_WB_RegBank_12_2_port, 
      pipeline_RegFile_DEC_WB_RegBank_12_3_port, 
      pipeline_RegFile_DEC_WB_RegBank_12_4_port, 
      pipeline_RegFile_DEC_WB_RegBank_12_5_port, 
      pipeline_RegFile_DEC_WB_RegBank_12_6_port, 
      pipeline_RegFile_DEC_WB_RegBank_12_7_port, 
      pipeline_RegFile_DEC_WB_RegBank_12_8_port, 
      pipeline_RegFile_DEC_WB_RegBank_12_9_port, 
      pipeline_RegFile_DEC_WB_RegBank_12_10_port, 
      pipeline_RegFile_DEC_WB_RegBank_12_11_port, 
      pipeline_RegFile_DEC_WB_RegBank_12_12_port, 
      pipeline_RegFile_DEC_WB_RegBank_12_13_port, 
      pipeline_RegFile_DEC_WB_RegBank_12_14_port, 
      pipeline_RegFile_DEC_WB_RegBank_12_15_port, 
      pipeline_RegFile_DEC_WB_RegBank_12_16_port, 
      pipeline_RegFile_DEC_WB_RegBank_12_17_port, 
      pipeline_RegFile_DEC_WB_RegBank_12_18_port, 
      pipeline_RegFile_DEC_WB_RegBank_12_19_port, 
      pipeline_RegFile_DEC_WB_RegBank_12_20_port, 
      pipeline_RegFile_DEC_WB_RegBank_12_21_port, 
      pipeline_RegFile_DEC_WB_RegBank_12_22_port, 
      pipeline_RegFile_DEC_WB_RegBank_12_23_port, 
      pipeline_RegFile_DEC_WB_RegBank_12_24_port, 
      pipeline_RegFile_DEC_WB_RegBank_12_25_port, 
      pipeline_RegFile_DEC_WB_RegBank_12_26_port, 
      pipeline_RegFile_DEC_WB_RegBank_12_27_port, 
      pipeline_RegFile_DEC_WB_RegBank_12_28_port, 
      pipeline_RegFile_DEC_WB_RegBank_12_29_port, 
      pipeline_RegFile_DEC_WB_RegBank_12_30_port, 
      pipeline_RegFile_DEC_WB_RegBank_12_31_port, 
      pipeline_RegFile_DEC_WB_RegBank_11_0_port, 
      pipeline_RegFile_DEC_WB_RegBank_11_1_port, 
      pipeline_RegFile_DEC_WB_RegBank_11_2_port, 
      pipeline_RegFile_DEC_WB_RegBank_11_3_port, 
      pipeline_RegFile_DEC_WB_RegBank_11_4_port, 
      pipeline_RegFile_DEC_WB_RegBank_11_5_port, 
      pipeline_RegFile_DEC_WB_RegBank_11_6_port, 
      pipeline_RegFile_DEC_WB_RegBank_11_7_port, 
      pipeline_RegFile_DEC_WB_RegBank_11_8_port, 
      pipeline_RegFile_DEC_WB_RegBank_11_9_port, 
      pipeline_RegFile_DEC_WB_RegBank_11_10_port, 
      pipeline_RegFile_DEC_WB_RegBank_11_11_port, 
      pipeline_RegFile_DEC_WB_RegBank_11_12_port, 
      pipeline_RegFile_DEC_WB_RegBank_11_13_port, 
      pipeline_RegFile_DEC_WB_RegBank_11_14_port, 
      pipeline_RegFile_DEC_WB_RegBank_11_15_port, 
      pipeline_RegFile_DEC_WB_RegBank_11_16_port, 
      pipeline_RegFile_DEC_WB_RegBank_11_17_port, 
      pipeline_RegFile_DEC_WB_RegBank_11_18_port, 
      pipeline_RegFile_DEC_WB_RegBank_11_19_port, 
      pipeline_RegFile_DEC_WB_RegBank_11_20_port, 
      pipeline_RegFile_DEC_WB_RegBank_11_21_port, 
      pipeline_RegFile_DEC_WB_RegBank_11_22_port, 
      pipeline_RegFile_DEC_WB_RegBank_11_23_port, 
      pipeline_RegFile_DEC_WB_RegBank_11_24_port, 
      pipeline_RegFile_DEC_WB_RegBank_11_25_port, 
      pipeline_RegFile_DEC_WB_RegBank_11_26_port, 
      pipeline_RegFile_DEC_WB_RegBank_11_27_port, 
      pipeline_RegFile_DEC_WB_RegBank_11_28_port, 
      pipeline_RegFile_DEC_WB_RegBank_11_29_port, 
      pipeline_RegFile_DEC_WB_RegBank_11_30_port, 
      pipeline_RegFile_DEC_WB_RegBank_11_31_port, 
      pipeline_RegFile_DEC_WB_RegBank_10_0_port, 
      pipeline_RegFile_DEC_WB_RegBank_10_1_port, 
      pipeline_RegFile_DEC_WB_RegBank_10_2_port, 
      pipeline_RegFile_DEC_WB_RegBank_10_3_port, 
      pipeline_RegFile_DEC_WB_RegBank_10_4_port, 
      pipeline_RegFile_DEC_WB_RegBank_10_5_port, 
      pipeline_RegFile_DEC_WB_RegBank_10_6_port, 
      pipeline_RegFile_DEC_WB_RegBank_10_7_port, 
      pipeline_RegFile_DEC_WB_RegBank_10_8_port, 
      pipeline_RegFile_DEC_WB_RegBank_10_9_port, 
      pipeline_RegFile_DEC_WB_RegBank_10_10_port, 
      pipeline_RegFile_DEC_WB_RegBank_10_11_port, 
      pipeline_RegFile_DEC_WB_RegBank_10_12_port, 
      pipeline_RegFile_DEC_WB_RegBank_10_13_port, 
      pipeline_RegFile_DEC_WB_RegBank_10_14_port, 
      pipeline_RegFile_DEC_WB_RegBank_10_15_port, 
      pipeline_RegFile_DEC_WB_RegBank_10_16_port, 
      pipeline_RegFile_DEC_WB_RegBank_10_17_port, 
      pipeline_RegFile_DEC_WB_RegBank_10_18_port, 
      pipeline_RegFile_DEC_WB_RegBank_10_19_port, 
      pipeline_RegFile_DEC_WB_RegBank_10_20_port, 
      pipeline_RegFile_DEC_WB_RegBank_10_21_port, 
      pipeline_RegFile_DEC_WB_RegBank_10_22_port, 
      pipeline_RegFile_DEC_WB_RegBank_10_23_port, 
      pipeline_RegFile_DEC_WB_RegBank_10_24_port, 
      pipeline_RegFile_DEC_WB_RegBank_10_25_port, 
      pipeline_RegFile_DEC_WB_RegBank_10_26_port, 
      pipeline_RegFile_DEC_WB_RegBank_10_27_port, 
      pipeline_RegFile_DEC_WB_RegBank_10_28_port, 
      pipeline_RegFile_DEC_WB_RegBank_10_29_port, 
      pipeline_RegFile_DEC_WB_RegBank_10_30_port, 
      pipeline_RegFile_DEC_WB_RegBank_10_31_port, 
      pipeline_RegFile_DEC_WB_RegBank_9_0_port, 
      pipeline_RegFile_DEC_WB_RegBank_9_1_port, 
      pipeline_RegFile_DEC_WB_RegBank_9_2_port, 
      pipeline_RegFile_DEC_WB_RegBank_9_3_port, 
      pipeline_RegFile_DEC_WB_RegBank_9_4_port, 
      pipeline_RegFile_DEC_WB_RegBank_9_5_port, 
      pipeline_RegFile_DEC_WB_RegBank_9_6_port, 
      pipeline_RegFile_DEC_WB_RegBank_9_7_port, 
      pipeline_RegFile_DEC_WB_RegBank_9_8_port, 
      pipeline_RegFile_DEC_WB_RegBank_9_9_port, 
      pipeline_RegFile_DEC_WB_RegBank_9_10_port, 
      pipeline_RegFile_DEC_WB_RegBank_9_11_port, 
      pipeline_RegFile_DEC_WB_RegBank_9_12_port, 
      pipeline_RegFile_DEC_WB_RegBank_9_13_port, 
      pipeline_RegFile_DEC_WB_RegBank_9_14_port, 
      pipeline_RegFile_DEC_WB_RegBank_9_15_port, 
      pipeline_RegFile_DEC_WB_RegBank_9_16_port, 
      pipeline_RegFile_DEC_WB_RegBank_9_17_port, 
      pipeline_RegFile_DEC_WB_RegBank_9_18_port, 
      pipeline_RegFile_DEC_WB_RegBank_9_19_port, 
      pipeline_RegFile_DEC_WB_RegBank_9_20_port, 
      pipeline_RegFile_DEC_WB_RegBank_9_21_port, 
      pipeline_RegFile_DEC_WB_RegBank_9_22_port, 
      pipeline_RegFile_DEC_WB_RegBank_9_23_port, 
      pipeline_RegFile_DEC_WB_RegBank_9_24_port, 
      pipeline_RegFile_DEC_WB_RegBank_9_25_port, 
      pipeline_RegFile_DEC_WB_RegBank_9_26_port, 
      pipeline_RegFile_DEC_WB_RegBank_9_27_port, 
      pipeline_RegFile_DEC_WB_RegBank_9_28_port, 
      pipeline_RegFile_DEC_WB_RegBank_9_29_port, 
      pipeline_RegFile_DEC_WB_RegBank_9_30_port, 
      pipeline_RegFile_DEC_WB_RegBank_9_31_port, 
      pipeline_RegFile_DEC_WB_RegBank_8_0_port, 
      pipeline_RegFile_DEC_WB_RegBank_8_1_port, 
      pipeline_RegFile_DEC_WB_RegBank_8_2_port, 
      pipeline_RegFile_DEC_WB_RegBank_8_3_port, 
      pipeline_RegFile_DEC_WB_RegBank_8_4_port, 
      pipeline_RegFile_DEC_WB_RegBank_8_5_port, 
      pipeline_RegFile_DEC_WB_RegBank_8_6_port, 
      pipeline_RegFile_DEC_WB_RegBank_8_7_port, 
      pipeline_RegFile_DEC_WB_RegBank_8_8_port, 
      pipeline_RegFile_DEC_WB_RegBank_8_9_port, 
      pipeline_RegFile_DEC_WB_RegBank_8_10_port, 
      pipeline_RegFile_DEC_WB_RegBank_8_11_port, 
      pipeline_RegFile_DEC_WB_RegBank_8_12_port, 
      pipeline_RegFile_DEC_WB_RegBank_8_13_port, 
      pipeline_RegFile_DEC_WB_RegBank_8_14_port, 
      pipeline_RegFile_DEC_WB_RegBank_8_15_port, 
      pipeline_RegFile_DEC_WB_RegBank_8_16_port, 
      pipeline_RegFile_DEC_WB_RegBank_8_17_port, 
      pipeline_RegFile_DEC_WB_RegBank_8_18_port, 
      pipeline_RegFile_DEC_WB_RegBank_8_19_port, 
      pipeline_RegFile_DEC_WB_RegBank_8_20_port, 
      pipeline_RegFile_DEC_WB_RegBank_8_21_port, 
      pipeline_RegFile_DEC_WB_RegBank_8_22_port, 
      pipeline_RegFile_DEC_WB_RegBank_8_23_port, 
      pipeline_RegFile_DEC_WB_RegBank_8_24_port, 
      pipeline_RegFile_DEC_WB_RegBank_8_25_port, 
      pipeline_RegFile_DEC_WB_RegBank_8_26_port, 
      pipeline_RegFile_DEC_WB_RegBank_8_27_port, 
      pipeline_RegFile_DEC_WB_RegBank_8_28_port, 
      pipeline_RegFile_DEC_WB_RegBank_8_29_port, 
      pipeline_RegFile_DEC_WB_RegBank_8_30_port, 
      pipeline_RegFile_DEC_WB_RegBank_8_31_port, 
      pipeline_RegFile_DEC_WB_RegBank_7_0_port, 
      pipeline_RegFile_DEC_WB_RegBank_7_1_port, 
      pipeline_RegFile_DEC_WB_RegBank_7_2_port, 
      pipeline_RegFile_DEC_WB_RegBank_7_3_port, 
      pipeline_RegFile_DEC_WB_RegBank_7_4_port, 
      pipeline_RegFile_DEC_WB_RegBank_7_5_port, 
      pipeline_RegFile_DEC_WB_RegBank_7_6_port, 
      pipeline_RegFile_DEC_WB_RegBank_7_7_port, 
      pipeline_RegFile_DEC_WB_RegBank_7_8_port, 
      pipeline_RegFile_DEC_WB_RegBank_7_9_port, 
      pipeline_RegFile_DEC_WB_RegBank_7_10_port, 
      pipeline_RegFile_DEC_WB_RegBank_7_11_port, 
      pipeline_RegFile_DEC_WB_RegBank_7_12_port, 
      pipeline_RegFile_DEC_WB_RegBank_7_13_port, 
      pipeline_RegFile_DEC_WB_RegBank_7_14_port, 
      pipeline_RegFile_DEC_WB_RegBank_7_15_port, 
      pipeline_RegFile_DEC_WB_RegBank_7_16_port, 
      pipeline_RegFile_DEC_WB_RegBank_7_17_port, 
      pipeline_RegFile_DEC_WB_RegBank_7_18_port, 
      pipeline_RegFile_DEC_WB_RegBank_7_19_port, 
      pipeline_RegFile_DEC_WB_RegBank_7_20_port, 
      pipeline_RegFile_DEC_WB_RegBank_7_21_port, 
      pipeline_RegFile_DEC_WB_RegBank_7_22_port, 
      pipeline_RegFile_DEC_WB_RegBank_7_23_port, 
      pipeline_RegFile_DEC_WB_RegBank_7_24_port, 
      pipeline_RegFile_DEC_WB_RegBank_7_25_port, 
      pipeline_RegFile_DEC_WB_RegBank_7_26_port, 
      pipeline_RegFile_DEC_WB_RegBank_7_27_port, 
      pipeline_RegFile_DEC_WB_RegBank_7_28_port, 
      pipeline_RegFile_DEC_WB_RegBank_7_29_port, 
      pipeline_RegFile_DEC_WB_RegBank_7_30_port, 
      pipeline_RegFile_DEC_WB_RegBank_7_31_port, 
      pipeline_RegFile_DEC_WB_RegBank_6_0_port, 
      pipeline_RegFile_DEC_WB_RegBank_6_1_port, 
      pipeline_RegFile_DEC_WB_RegBank_6_2_port, 
      pipeline_RegFile_DEC_WB_RegBank_6_3_port, 
      pipeline_RegFile_DEC_WB_RegBank_6_4_port, 
      pipeline_RegFile_DEC_WB_RegBank_6_5_port, 
      pipeline_RegFile_DEC_WB_RegBank_6_6_port, 
      pipeline_RegFile_DEC_WB_RegBank_6_7_port, 
      pipeline_RegFile_DEC_WB_RegBank_6_8_port, 
      pipeline_RegFile_DEC_WB_RegBank_6_9_port, 
      pipeline_RegFile_DEC_WB_RegBank_6_10_port, 
      pipeline_RegFile_DEC_WB_RegBank_6_11_port, 
      pipeline_RegFile_DEC_WB_RegBank_6_12_port, 
      pipeline_RegFile_DEC_WB_RegBank_6_13_port, 
      pipeline_RegFile_DEC_WB_RegBank_6_14_port, 
      pipeline_RegFile_DEC_WB_RegBank_6_15_port, 
      pipeline_RegFile_DEC_WB_RegBank_6_16_port, 
      pipeline_RegFile_DEC_WB_RegBank_6_17_port, 
      pipeline_RegFile_DEC_WB_RegBank_6_18_port, 
      pipeline_RegFile_DEC_WB_RegBank_6_19_port, 
      pipeline_RegFile_DEC_WB_RegBank_6_20_port, 
      pipeline_RegFile_DEC_WB_RegBank_6_21_port, 
      pipeline_RegFile_DEC_WB_RegBank_6_22_port, 
      pipeline_RegFile_DEC_WB_RegBank_6_23_port, 
      pipeline_RegFile_DEC_WB_RegBank_6_24_port, 
      pipeline_RegFile_DEC_WB_RegBank_6_25_port, 
      pipeline_RegFile_DEC_WB_RegBank_6_26_port, 
      pipeline_RegFile_DEC_WB_RegBank_6_27_port, 
      pipeline_RegFile_DEC_WB_RegBank_6_28_port, 
      pipeline_RegFile_DEC_WB_RegBank_6_29_port, 
      pipeline_RegFile_DEC_WB_RegBank_6_30_port, 
      pipeline_RegFile_DEC_WB_RegBank_6_31_port, 
      pipeline_RegFile_DEC_WB_RegBank_5_0_port, 
      pipeline_RegFile_DEC_WB_RegBank_5_1_port, 
      pipeline_RegFile_DEC_WB_RegBank_5_2_port, 
      pipeline_RegFile_DEC_WB_RegBank_5_3_port, 
      pipeline_RegFile_DEC_WB_RegBank_5_4_port, 
      pipeline_RegFile_DEC_WB_RegBank_5_5_port, 
      pipeline_RegFile_DEC_WB_RegBank_5_6_port, 
      pipeline_RegFile_DEC_WB_RegBank_5_7_port, 
      pipeline_RegFile_DEC_WB_RegBank_5_8_port, 
      pipeline_RegFile_DEC_WB_RegBank_5_9_port, 
      pipeline_RegFile_DEC_WB_RegBank_5_10_port, 
      pipeline_RegFile_DEC_WB_RegBank_5_11_port, 
      pipeline_RegFile_DEC_WB_RegBank_5_12_port, 
      pipeline_RegFile_DEC_WB_RegBank_5_13_port, 
      pipeline_RegFile_DEC_WB_RegBank_5_14_port, 
      pipeline_RegFile_DEC_WB_RegBank_5_15_port, 
      pipeline_RegFile_DEC_WB_RegBank_5_16_port, 
      pipeline_RegFile_DEC_WB_RegBank_5_17_port, 
      pipeline_RegFile_DEC_WB_RegBank_5_18_port, 
      pipeline_RegFile_DEC_WB_RegBank_5_19_port, 
      pipeline_RegFile_DEC_WB_RegBank_5_20_port, 
      pipeline_RegFile_DEC_WB_RegBank_5_21_port, 
      pipeline_RegFile_DEC_WB_RegBank_5_22_port, 
      pipeline_RegFile_DEC_WB_RegBank_5_23_port, 
      pipeline_RegFile_DEC_WB_RegBank_5_24_port, 
      pipeline_RegFile_DEC_WB_RegBank_5_25_port, 
      pipeline_RegFile_DEC_WB_RegBank_5_26_port, 
      pipeline_RegFile_DEC_WB_RegBank_5_27_port, 
      pipeline_RegFile_DEC_WB_RegBank_5_28_port, 
      pipeline_RegFile_DEC_WB_RegBank_5_29_port, 
      pipeline_RegFile_DEC_WB_RegBank_5_30_port, 
      pipeline_RegFile_DEC_WB_RegBank_5_31_port, 
      pipeline_RegFile_DEC_WB_RegBank_4_0_port, 
      pipeline_RegFile_DEC_WB_RegBank_4_1_port, 
      pipeline_RegFile_DEC_WB_RegBank_4_2_port, 
      pipeline_RegFile_DEC_WB_RegBank_4_3_port, 
      pipeline_RegFile_DEC_WB_RegBank_4_4_port, 
      pipeline_RegFile_DEC_WB_RegBank_4_5_port, 
      pipeline_RegFile_DEC_WB_RegBank_4_6_port, 
      pipeline_RegFile_DEC_WB_RegBank_4_7_port, 
      pipeline_RegFile_DEC_WB_RegBank_4_8_port, 
      pipeline_RegFile_DEC_WB_RegBank_4_9_port, 
      pipeline_RegFile_DEC_WB_RegBank_4_10_port, 
      pipeline_RegFile_DEC_WB_RegBank_4_11_port, 
      pipeline_RegFile_DEC_WB_RegBank_4_12_port, 
      pipeline_RegFile_DEC_WB_RegBank_4_13_port, 
      pipeline_RegFile_DEC_WB_RegBank_4_14_port, 
      pipeline_RegFile_DEC_WB_RegBank_4_15_port, 
      pipeline_RegFile_DEC_WB_RegBank_4_16_port, 
      pipeline_RegFile_DEC_WB_RegBank_4_17_port, 
      pipeline_RegFile_DEC_WB_RegBank_4_18_port, 
      pipeline_RegFile_DEC_WB_RegBank_4_19_port, 
      pipeline_RegFile_DEC_WB_RegBank_4_20_port, 
      pipeline_RegFile_DEC_WB_RegBank_4_21_port, 
      pipeline_RegFile_DEC_WB_RegBank_4_22_port, 
      pipeline_RegFile_DEC_WB_RegBank_4_23_port, 
      pipeline_RegFile_DEC_WB_RegBank_4_24_port, 
      pipeline_RegFile_DEC_WB_RegBank_4_25_port, 
      pipeline_RegFile_DEC_WB_RegBank_4_26_port, 
      pipeline_RegFile_DEC_WB_RegBank_4_27_port, 
      pipeline_RegFile_DEC_WB_RegBank_4_28_port, 
      pipeline_RegFile_DEC_WB_RegBank_4_29_port, 
      pipeline_RegFile_DEC_WB_RegBank_4_30_port, 
      pipeline_RegFile_DEC_WB_RegBank_4_31_port, 
      pipeline_RegFile_DEC_WB_RegBank_3_0_port, 
      pipeline_RegFile_DEC_WB_RegBank_3_1_port, 
      pipeline_RegFile_DEC_WB_RegBank_3_2_port, 
      pipeline_RegFile_DEC_WB_RegBank_3_3_port, 
      pipeline_RegFile_DEC_WB_RegBank_3_4_port, 
      pipeline_RegFile_DEC_WB_RegBank_3_5_port, 
      pipeline_RegFile_DEC_WB_RegBank_3_6_port, 
      pipeline_RegFile_DEC_WB_RegBank_3_7_port, 
      pipeline_RegFile_DEC_WB_RegBank_3_8_port, 
      pipeline_RegFile_DEC_WB_RegBank_3_9_port, 
      pipeline_RegFile_DEC_WB_RegBank_3_10_port, 
      pipeline_RegFile_DEC_WB_RegBank_3_11_port, 
      pipeline_RegFile_DEC_WB_RegBank_3_12_port, 
      pipeline_RegFile_DEC_WB_RegBank_3_13_port, 
      pipeline_RegFile_DEC_WB_RegBank_3_14_port, 
      pipeline_RegFile_DEC_WB_RegBank_3_15_port, 
      pipeline_RegFile_DEC_WB_RegBank_3_16_port, 
      pipeline_RegFile_DEC_WB_RegBank_3_17_port, 
      pipeline_RegFile_DEC_WB_RegBank_3_18_port, 
      pipeline_RegFile_DEC_WB_RegBank_3_19_port, 
      pipeline_RegFile_DEC_WB_RegBank_3_20_port, 
      pipeline_RegFile_DEC_WB_RegBank_3_21_port, 
      pipeline_RegFile_DEC_WB_RegBank_3_22_port, 
      pipeline_RegFile_DEC_WB_RegBank_3_23_port, 
      pipeline_RegFile_DEC_WB_RegBank_3_24_port, 
      pipeline_RegFile_DEC_WB_RegBank_3_25_port, 
      pipeline_RegFile_DEC_WB_RegBank_3_26_port, 
      pipeline_RegFile_DEC_WB_RegBank_3_27_port, 
      pipeline_RegFile_DEC_WB_RegBank_3_28_port, 
      pipeline_RegFile_DEC_WB_RegBank_3_29_port, 
      pipeline_RegFile_DEC_WB_RegBank_3_30_port, 
      pipeline_RegFile_DEC_WB_RegBank_3_31_port, 
      pipeline_RegFile_DEC_WB_RegBank_2_0_port, 
      pipeline_RegFile_DEC_WB_RegBank_2_1_port, 
      pipeline_RegFile_DEC_WB_RegBank_2_2_port, 
      pipeline_RegFile_DEC_WB_RegBank_2_3_port, 
      pipeline_RegFile_DEC_WB_RegBank_2_4_port, 
      pipeline_RegFile_DEC_WB_RegBank_2_5_port, 
      pipeline_RegFile_DEC_WB_RegBank_2_6_port, 
      pipeline_RegFile_DEC_WB_RegBank_2_7_port, 
      pipeline_RegFile_DEC_WB_RegBank_2_8_port, 
      pipeline_RegFile_DEC_WB_RegBank_2_9_port, 
      pipeline_RegFile_DEC_WB_RegBank_2_10_port, 
      pipeline_RegFile_DEC_WB_RegBank_2_11_port, 
      pipeline_RegFile_DEC_WB_RegBank_2_12_port, 
      pipeline_RegFile_DEC_WB_RegBank_2_13_port, 
      pipeline_RegFile_DEC_WB_RegBank_2_14_port, 
      pipeline_RegFile_DEC_WB_RegBank_2_15_port, 
      pipeline_RegFile_DEC_WB_RegBank_2_16_port, 
      pipeline_RegFile_DEC_WB_RegBank_2_17_port, 
      pipeline_RegFile_DEC_WB_RegBank_2_18_port, 
      pipeline_RegFile_DEC_WB_RegBank_2_19_port, 
      pipeline_RegFile_DEC_WB_RegBank_2_20_port, 
      pipeline_RegFile_DEC_WB_RegBank_2_21_port, 
      pipeline_RegFile_DEC_WB_RegBank_2_22_port, 
      pipeline_RegFile_DEC_WB_RegBank_2_23_port, 
      pipeline_RegFile_DEC_WB_RegBank_2_24_port, 
      pipeline_RegFile_DEC_WB_RegBank_2_25_port, 
      pipeline_RegFile_DEC_WB_RegBank_2_26_port, 
      pipeline_RegFile_DEC_WB_RegBank_2_27_port, 
      pipeline_RegFile_DEC_WB_RegBank_2_28_port, 
      pipeline_RegFile_DEC_WB_RegBank_2_29_port, 
      pipeline_RegFile_DEC_WB_RegBank_2_30_port, 
      pipeline_RegFile_DEC_WB_RegBank_2_31_port, 
      pipeline_RegFile_DEC_WB_RegBank_1_0_port, 
      pipeline_RegFile_DEC_WB_RegBank_1_1_port, 
      pipeline_RegFile_DEC_WB_RegBank_1_2_port, 
      pipeline_RegFile_DEC_WB_RegBank_1_3_port, 
      pipeline_RegFile_DEC_WB_RegBank_1_4_port, 
      pipeline_RegFile_DEC_WB_RegBank_1_5_port, 
      pipeline_RegFile_DEC_WB_RegBank_1_6_port, 
      pipeline_RegFile_DEC_WB_RegBank_1_7_port, 
      pipeline_RegFile_DEC_WB_RegBank_1_8_port, 
      pipeline_RegFile_DEC_WB_RegBank_1_9_port, 
      pipeline_RegFile_DEC_WB_RegBank_1_10_port, 
      pipeline_RegFile_DEC_WB_RegBank_1_11_port, 
      pipeline_RegFile_DEC_WB_RegBank_1_12_port, 
      pipeline_RegFile_DEC_WB_RegBank_1_13_port, 
      pipeline_RegFile_DEC_WB_RegBank_1_14_port, 
      pipeline_RegFile_DEC_WB_RegBank_1_15_port, 
      pipeline_RegFile_DEC_WB_RegBank_1_16_port, 
      pipeline_RegFile_DEC_WB_RegBank_1_17_port, 
      pipeline_RegFile_DEC_WB_RegBank_1_18_port, 
      pipeline_RegFile_DEC_WB_RegBank_1_19_port, 
      pipeline_RegFile_DEC_WB_RegBank_1_20_port, 
      pipeline_RegFile_DEC_WB_RegBank_1_21_port, 
      pipeline_RegFile_DEC_WB_RegBank_1_22_port, 
      pipeline_RegFile_DEC_WB_RegBank_1_23_port, 
      pipeline_RegFile_DEC_WB_RegBank_1_24_port, 
      pipeline_RegFile_DEC_WB_RegBank_1_25_port, 
      pipeline_RegFile_DEC_WB_RegBank_1_26_port, 
      pipeline_RegFile_DEC_WB_RegBank_1_27_port, 
      pipeline_RegFile_DEC_WB_RegBank_1_28_port, 
      pipeline_RegFile_DEC_WB_RegBank_1_29_port, 
      pipeline_RegFile_DEC_WB_RegBank_1_30_port, 
      pipeline_RegFile_DEC_WB_RegBank_1_31_port, pipeline_IDEX_Stage_N217, 
      pipeline_IDEX_Stage_N216, pipeline_IDEX_Stage_N215, 
      pipeline_IDEX_Stage_N214, pipeline_IDEX_Stage_N213, 
      pipeline_IDEX_Stage_N212, pipeline_IDEX_Stage_N211, 
      pipeline_IDEX_Stage_N210, pipeline_IDEX_Stage_N209, 
      pipeline_IDEX_Stage_N208, pipeline_IDEX_Stage_N207, 
      pipeline_IDEX_Stage_N206, pipeline_IDEX_Stage_N205, 
      pipeline_IDEX_Stage_N204, pipeline_IDEX_Stage_N203, 
      pipeline_IDEX_Stage_N202, pipeline_IDEX_Stage_N201, 
      pipeline_IDEX_Stage_N200, pipeline_IDEX_Stage_N199, 
      pipeline_IDEX_Stage_N198, pipeline_IDEX_Stage_N197, 
      pipeline_IDEX_Stage_N181, pipeline_IDEX_Stage_N180, 
      pipeline_IDEX_Stage_N179, pipeline_IDEX_Stage_N178, 
      pipeline_IDEX_Stage_N177, pipeline_IDEX_Stage_N176, 
      pipeline_IDEX_Stage_N175, pipeline_IDEX_Stage_N174, 
      pipeline_IDEX_Stage_N173, pipeline_IDEX_Stage_N172, 
      pipeline_IDEX_Stage_N171, pipeline_IDEX_Stage_N170, 
      pipeline_IDEX_Stage_N169, pipeline_IDEX_Stage_N168, 
      pipeline_IDEX_Stage_N167, pipeline_IDEX_Stage_N166, 
      pipeline_IDEX_Stage_N165, pipeline_IDEX_Stage_N164, 
      pipeline_IDEX_Stage_N163, pipeline_IDEX_Stage_N162, 
      pipeline_IDEX_Stage_N161, pipeline_IDEX_Stage_N160, 
      pipeline_IDEX_Stage_N159, pipeline_IDEX_Stage_N158, 
      pipeline_IDEX_Stage_N157, pipeline_IDEX_Stage_N156, 
      pipeline_IDEX_Stage_N155, pipeline_IDEX_Stage_N154, 
      pipeline_IDEX_Stage_N153, pipeline_IDEX_Stage_N152, 
      pipeline_IDEX_Stage_N151, pipeline_IDEX_Stage_N150, 
      pipeline_IDEX_Stage_N149, pipeline_IDEX_Stage_N148, 
      pipeline_IDEX_Stage_N147, pipeline_IDEX_Stage_N146, 
      pipeline_IDEX_Stage_N145, pipeline_IDEX_Stage_N144, 
      pipeline_IDEX_Stage_N143, pipeline_IDEX_Stage_N142, 
      pipeline_IDEX_Stage_N141, pipeline_IDEX_Stage_N140, 
      pipeline_IDEX_Stage_N139, pipeline_IDEX_Stage_N138, 
      pipeline_IDEX_Stage_N137, pipeline_IDEX_Stage_N136, 
      pipeline_IDEX_Stage_N135, pipeline_IDEX_Stage_N134, 
      pipeline_IDEX_Stage_N133, pipeline_IDEX_Stage_N132, 
      pipeline_IDEX_Stage_N131, pipeline_IDEX_Stage_N130, 
      pipeline_IDEX_Stage_N129, pipeline_IDEX_Stage_N128, 
      pipeline_IDEX_Stage_N127, pipeline_IDEX_Stage_N126, 
      pipeline_IDEX_Stage_N125, pipeline_IDEX_Stage_N124, 
      pipeline_IDEX_Stage_N123, pipeline_IDEX_Stage_N122, 
      pipeline_IDEX_Stage_N121, pipeline_IDEX_Stage_N120, 
      pipeline_IDEX_Stage_N119, pipeline_IDEX_Stage_N118, 
      pipeline_IDEX_Stage_N117, pipeline_IDEX_Stage_N116, 
      pipeline_IDEX_Stage_N115, pipeline_IDEX_Stage_N114, 
      pipeline_IDEX_Stage_N113, pipeline_IDEX_Stage_N112, 
      pipeline_IDEX_Stage_N111, pipeline_IDEX_Stage_N110, 
      pipeline_IDEX_Stage_N109, pipeline_IDEX_Stage_N108, 
      pipeline_IDEX_Stage_N107, pipeline_IDEX_Stage_N106, 
      pipeline_IDEX_Stage_N105, pipeline_IDEX_Stage_N104, 
      pipeline_IDEX_Stage_N103, pipeline_IDEX_Stage_N102, 
      pipeline_IDEX_Stage_N101, pipeline_IDEX_Stage_N100, 
      pipeline_IDEX_Stage_N99, pipeline_IDEX_Stage_N98, pipeline_IDEX_Stage_N97
      , pipeline_IDEX_Stage_N96, pipeline_IDEX_Stage_N95, 
      pipeline_IDEX_Stage_N94, pipeline_IDEX_Stage_N93, pipeline_IDEX_Stage_N92
      , pipeline_IDEX_Stage_N91, pipeline_IDEX_Stage_N90, 
      pipeline_IDEX_Stage_N89, pipeline_stageE_input2_to_ALU_0_port, 
      pipeline_stageE_input1_to_ALU_1_port, 
      pipeline_stageE_input1_to_ALU_3_port, 
      pipeline_stageE_input1_to_ALU_4_port, 
      pipeline_stageE_input1_to_ALU_5_port, 
      pipeline_stageE_input1_to_ALU_6_port, 
      pipeline_stageE_input1_to_ALU_7_port, 
      pipeline_stageE_input1_to_ALU_8_port, 
      pipeline_stageE_input1_to_ALU_9_port, 
      pipeline_stageE_input1_to_ALU_10_port, 
      pipeline_stageE_input1_to_ALU_11_port, 
      pipeline_stageE_input1_to_ALU_12_port, 
      pipeline_stageE_input1_to_ALU_13_port, 
      pipeline_stageE_input1_to_ALU_14_port, 
      pipeline_stageE_input1_to_ALU_15_port, 
      pipeline_stageE_input1_to_ALU_16_port, 
      pipeline_stageE_input1_to_ALU_17_port, 
      pipeline_stageE_input1_to_ALU_18_port, 
      pipeline_stageE_input1_to_ALU_19_port, 
      pipeline_stageE_input1_to_ALU_20_port, 
      pipeline_stageE_input1_to_ALU_21_port, 
      pipeline_stageE_input1_to_ALU_22_port, 
      pipeline_stageE_input1_to_ALU_23_port, 
      pipeline_stageE_input1_to_ALU_24_port, 
      pipeline_stageE_input1_to_ALU_25_port, 
      pipeline_stageE_input1_to_ALU_26_port, 
      pipeline_stageE_input1_to_ALU_27_port, 
      pipeline_stageE_input1_to_ALU_28_port, 
      pipeline_stageE_input1_to_ALU_29_port, 
      pipeline_stageE_input1_to_ALU_30_port, 
      pipeline_stageE_EXE_ALU_add_alu_sCout_0_port, 
      pipeline_stageE_EXE_ALU_alu_shift_N265, 
      pipeline_stageE_EXE_ALU_alu_shift_N264, 
      pipeline_stageE_EXE_ALU_alu_shift_N263, 
      pipeline_stageE_EXE_ALU_alu_shift_N262, 
      pipeline_stageE_EXE_ALU_alu_shift_N261, 
      pipeline_stageE_EXE_ALU_alu_shift_N260, 
      pipeline_stageE_EXE_ALU_alu_shift_N259, 
      pipeline_stageE_EXE_ALU_alu_shift_N258, 
      pipeline_stageE_EXE_ALU_alu_shift_N257, 
      pipeline_stageE_EXE_ALU_alu_shift_N256, 
      pipeline_stageE_EXE_ALU_alu_shift_N255, 
      pipeline_stageE_EXE_ALU_alu_shift_N254, 
      pipeline_stageE_EXE_ALU_alu_shift_N253, 
      pipeline_stageE_EXE_ALU_alu_shift_N252, 
      pipeline_stageE_EXE_ALU_alu_shift_N251, 
      pipeline_stageE_EXE_ALU_alu_shift_N250, 
      pipeline_stageE_EXE_ALU_alu_shift_N249, 
      pipeline_stageE_EXE_ALU_alu_shift_N248, 
      pipeline_stageE_EXE_ALU_alu_shift_N247, 
      pipeline_stageE_EXE_ALU_alu_shift_N246, 
      pipeline_stageE_EXE_ALU_alu_shift_N245, 
      pipeline_stageE_EXE_ALU_alu_shift_N244, 
      pipeline_stageE_EXE_ALU_alu_shift_N243, 
      pipeline_stageE_EXE_ALU_alu_shift_N242, 
      pipeline_stageE_EXE_ALU_alu_shift_N241, 
      pipeline_stageE_EXE_ALU_alu_shift_N240, 
      pipeline_stageE_EXE_ALU_alu_shift_N239, 
      pipeline_stageE_EXE_ALU_alu_shift_N238, 
      pipeline_stageE_EXE_ALU_alu_shift_N237, 
      pipeline_stageE_EXE_ALU_alu_shift_N236, 
      pipeline_stageE_EXE_ALU_alu_shift_N235, 
      pipeline_stageE_EXE_ALU_alu_shift_N234, 
      pipeline_stageE_EXE_ALU_alu_shift_N233, 
      pipeline_stageE_EXE_ALU_alu_shift_N232, 
      pipeline_stageE_EXE_ALU_alu_shift_N231, 
      pipeline_stageE_EXE_ALU_alu_shift_N230, 
      pipeline_stageE_EXE_ALU_alu_shift_N229, 
      pipeline_stageE_EXE_ALU_alu_shift_N228, 
      pipeline_stageE_EXE_ALU_alu_shift_N227, 
      pipeline_stageE_EXE_ALU_alu_shift_N226, 
      pipeline_stageE_EXE_ALU_alu_shift_N225, 
      pipeline_stageE_EXE_ALU_alu_shift_N224, 
      pipeline_stageE_EXE_ALU_alu_shift_N223, 
      pipeline_stageE_EXE_ALU_alu_shift_N222, 
      pipeline_stageE_EXE_ALU_alu_shift_N221, 
      pipeline_stageE_EXE_ALU_alu_shift_N220, 
      pipeline_stageE_EXE_ALU_alu_shift_N219, 
      pipeline_stageE_EXE_ALU_alu_shift_N218, 
      pipeline_stageE_EXE_ALU_alu_shift_N217, 
      pipeline_stageE_EXE_ALU_alu_shift_N216, 
      pipeline_stageE_EXE_ALU_alu_shift_N215, 
      pipeline_stageE_EXE_ALU_alu_shift_N214, 
      pipeline_stageE_EXE_ALU_alu_shift_N213, 
      pipeline_stageE_EXE_ALU_alu_shift_N212, 
      pipeline_stageE_EXE_ALU_alu_shift_N211, 
      pipeline_stageE_EXE_ALU_alu_shift_N210, 
      pipeline_stageE_EXE_ALU_alu_shift_N209, 
      pipeline_stageE_EXE_ALU_alu_shift_N208, 
      pipeline_stageE_EXE_ALU_alu_shift_N207, 
      pipeline_stageE_EXE_ALU_alu_shift_N206, 
      pipeline_stageE_EXE_ALU_alu_shift_N205, 
      pipeline_stageE_EXE_ALU_alu_shift_N204, 
      pipeline_stageE_EXE_ALU_alu_shift_N203, 
      pipeline_stageE_EXE_ALU_alu_shift_N202, 
      pipeline_stageE_EXE_ALU_alu_shift_N168, 
      pipeline_stageE_EXE_ALU_alu_shift_N167, 
      pipeline_stageE_EXE_ALU_alu_shift_N166, 
      pipeline_stageE_EXE_ALU_alu_shift_N165, 
      pipeline_stageE_EXE_ALU_alu_shift_N164, 
      pipeline_stageE_EXE_ALU_alu_shift_N163, 
      pipeline_stageE_EXE_ALU_alu_shift_N162, 
      pipeline_stageE_EXE_ALU_alu_shift_N161, 
      pipeline_stageE_EXE_ALU_alu_shift_N160, 
      pipeline_stageE_EXE_ALU_alu_shift_N159, 
      pipeline_stageE_EXE_ALU_alu_shift_N158, 
      pipeline_stageE_EXE_ALU_alu_shift_N157, 
      pipeline_stageE_EXE_ALU_alu_shift_N156, 
      pipeline_stageE_EXE_ALU_alu_shift_N155, 
      pipeline_stageE_EXE_ALU_alu_shift_N154, 
      pipeline_stageE_EXE_ALU_alu_shift_N153, 
      pipeline_stageE_EXE_ALU_alu_shift_N152, 
      pipeline_stageE_EXE_ALU_alu_shift_N151, 
      pipeline_stageE_EXE_ALU_alu_shift_N150, 
      pipeline_stageE_EXE_ALU_alu_shift_N149, 
      pipeline_stageE_EXE_ALU_alu_shift_N148, 
      pipeline_stageE_EXE_ALU_alu_shift_N147, 
      pipeline_stageE_EXE_ALU_alu_shift_N146, 
      pipeline_stageE_EXE_ALU_alu_shift_N145, 
      pipeline_stageE_EXE_ALU_alu_shift_N144, 
      pipeline_stageE_EXE_ALU_alu_shift_N143, 
      pipeline_stageE_EXE_ALU_alu_shift_N142, 
      pipeline_stageE_EXE_ALU_alu_shift_N141, 
      pipeline_stageE_EXE_ALU_alu_shift_N140, 
      pipeline_stageE_EXE_ALU_alu_shift_N139, 
      pipeline_stageE_EXE_ALU_alu_shift_N138, 
      pipeline_stageE_EXE_ALU_alu_shift_N137, 
      pipeline_stageE_EXE_ALU_alu_shift_N136, 
      pipeline_stageE_EXE_ALU_alu_shift_N135, 
      pipeline_stageE_EXE_ALU_alu_shift_N134, 
      pipeline_stageE_EXE_ALU_alu_shift_N133, 
      pipeline_stageE_EXE_ALU_alu_shift_N132, 
      pipeline_stageE_EXE_ALU_alu_shift_N131, 
      pipeline_stageE_EXE_ALU_alu_shift_N130, 
      pipeline_stageE_EXE_ALU_alu_shift_N129, 
      pipeline_stageE_EXE_ALU_alu_shift_N128, 
      pipeline_stageE_EXE_ALU_alu_shift_N127, 
      pipeline_stageE_EXE_ALU_alu_shift_N126, 
      pipeline_stageE_EXE_ALU_alu_shift_N125, 
      pipeline_stageE_EXE_ALU_alu_shift_N124, 
      pipeline_stageE_EXE_ALU_alu_shift_N123, 
      pipeline_stageE_EXE_ALU_alu_shift_N122, 
      pipeline_stageE_EXE_ALU_alu_shift_N121, 
      pipeline_stageE_EXE_ALU_alu_shift_N120, 
      pipeline_stageE_EXE_ALU_alu_shift_N119, 
      pipeline_stageE_EXE_ALU_alu_shift_N118, 
      pipeline_stageE_EXE_ALU_alu_shift_N117, 
      pipeline_stageE_EXE_ALU_alu_shift_N116, 
      pipeline_stageE_EXE_ALU_alu_shift_N115, 
      pipeline_stageE_EXE_ALU_alu_shift_N114, 
      pipeline_stageE_EXE_ALU_alu_shift_N113, 
      pipeline_stageE_EXE_ALU_alu_shift_N112, 
      pipeline_stageE_EXE_ALU_alu_shift_N111, 
      pipeline_stageE_EXE_ALU_alu_shift_N110, 
      pipeline_stageE_EXE_ALU_alu_shift_N109, 
      pipeline_stageE_EXE_ALU_alu_shift_N108, 
      pipeline_stageE_EXE_ALU_alu_shift_N107, 
      pipeline_stageE_EXE_ALU_alu_shift_N106, 
      pipeline_stageE_EXE_ALU_alu_shift_N105, 
      pipeline_stageE_EXE_ALU_alu_shift_N70, 
      pipeline_stageE_EXE_ALU_alu_shift_N69, 
      pipeline_stageE_EXE_ALU_alu_shift_N68, 
      pipeline_stageE_EXE_ALU_alu_shift_N67, 
      pipeline_stageE_EXE_ALU_alu_shift_N66, 
      pipeline_stageE_EXE_ALU_alu_shift_N65, 
      pipeline_stageE_EXE_ALU_alu_shift_N64, 
      pipeline_stageE_EXE_ALU_alu_shift_N63, 
      pipeline_stageE_EXE_ALU_alu_shift_N62, 
      pipeline_stageE_EXE_ALU_alu_shift_N61, 
      pipeline_stageE_EXE_ALU_alu_shift_N60, 
      pipeline_stageE_EXE_ALU_alu_shift_N59, 
      pipeline_stageE_EXE_ALU_alu_shift_N58, 
      pipeline_stageE_EXE_ALU_alu_shift_N57, 
      pipeline_stageE_EXE_ALU_alu_shift_N56, 
      pipeline_stageE_EXE_ALU_alu_shift_N55, 
      pipeline_stageE_EXE_ALU_alu_shift_N54, 
      pipeline_stageE_EXE_ALU_alu_shift_N53, 
      pipeline_stageE_EXE_ALU_alu_shift_N52, 
      pipeline_stageE_EXE_ALU_alu_shift_N51, 
      pipeline_stageE_EXE_ALU_alu_shift_N50, 
      pipeline_stageE_EXE_ALU_alu_shift_N49, 
      pipeline_stageE_EXE_ALU_alu_shift_N48, 
      pipeline_stageE_EXE_ALU_alu_shift_N47, 
      pipeline_stageE_EXE_ALU_alu_shift_N46, 
      pipeline_stageE_EXE_ALU_alu_shift_N45, 
      pipeline_stageE_EXE_ALU_alu_shift_N44, 
      pipeline_stageE_EXE_ALU_alu_shift_N43, 
      pipeline_stageE_EXE_ALU_alu_shift_N42, 
      pipeline_stageE_EXE_ALU_alu_shift_N41, 
      pipeline_stageE_EXE_ALU_alu_shift_N40, 
      pipeline_stageE_EXE_ALU_alu_shift_N39, 
      pipeline_stageE_EXE_ALU_alu_shift_N38, 
      pipeline_stageE_EXE_ALU_alu_shift_N37, 
      pipeline_stageE_EXE_ALU_alu_shift_N36, 
      pipeline_stageE_EXE_ALU_alu_shift_N35, 
      pipeline_stageE_EXE_ALU_alu_shift_N34, 
      pipeline_stageE_EXE_ALU_alu_shift_N33, 
      pipeline_stageE_EXE_ALU_alu_shift_N32, 
      pipeline_stageE_EXE_ALU_alu_shift_N31, 
      pipeline_stageE_EXE_ALU_alu_shift_N30, 
      pipeline_stageE_EXE_ALU_alu_shift_N29, 
      pipeline_stageE_EXE_ALU_alu_shift_N28, 
      pipeline_stageE_EXE_ALU_alu_shift_N27, 
      pipeline_stageE_EXE_ALU_alu_shift_N26, 
      pipeline_stageE_EXE_ALU_alu_shift_N25, 
      pipeline_stageE_EXE_ALU_alu_shift_N24, 
      pipeline_stageE_EXE_ALU_alu_shift_N23, 
      pipeline_stageE_EXE_ALU_alu_shift_N22, 
      pipeline_stageE_EXE_ALU_alu_shift_N21, 
      pipeline_stageE_EXE_ALU_alu_shift_N20, 
      pipeline_stageE_EXE_ALU_alu_shift_N19, 
      pipeline_stageE_EXE_ALU_alu_shift_N18, 
      pipeline_stageE_EXE_ALU_alu_shift_N17, 
      pipeline_stageE_EXE_ALU_alu_shift_N16, 
      pipeline_stageE_EXE_ALU_alu_shift_N15, 
      pipeline_stageE_EXE_ALU_alu_shift_N14, 
      pipeline_stageE_EXE_ALU_alu_shift_N13, 
      pipeline_stageE_EXE_ALU_alu_shift_N12, 
      pipeline_stageE_EXE_ALU_alu_shift_N11, 
      pipeline_stageE_EXE_ALU_alu_shift_N10, 
      pipeline_stageE_EXE_ALU_alu_shift_N9, 
      pipeline_stageE_EXE_ALU_alu_shift_N8, 
      pipeline_stageE_EXE_ALU_alu_shift_N7, pipeline_EXMEM_stage_N76, 
      pipeline_EXMEM_stage_N75, pipeline_EXMEM_stage_N74, 
      pipeline_EXMEM_stage_N73, pipeline_EXMEM_stage_N72, 
      pipeline_EXMEM_stage_N71, pipeline_EXMEM_stage_N70, 
      pipeline_EXMEM_stage_N69, pipeline_EXMEM_stage_N68, 
      pipeline_EXMEM_stage_N67, pipeline_EXMEM_stage_N66, 
      pipeline_EXMEM_stage_N65, pipeline_EXMEM_stage_N64, 
      pipeline_EXMEM_stage_N63, pipeline_EXMEM_stage_N62, 
      pipeline_EXMEM_stage_N61, pipeline_EXMEM_stage_N60, 
      pipeline_EXMEM_stage_N59, pipeline_EXMEM_stage_N58, 
      pipeline_EXMEM_stage_N57, pipeline_EXMEM_stage_N56, 
      pipeline_EXMEM_stage_N55, pipeline_EXMEM_stage_N54, 
      pipeline_EXMEM_stage_N53, pipeline_EXMEM_stage_N52, 
      pipeline_EXMEM_stage_N51, pipeline_EXMEM_stage_N50, 
      pipeline_EXMEM_stage_N49, pipeline_EXMEM_stage_N48, 
      pipeline_EXMEM_stage_N47, pipeline_EXMEM_stage_N46, 
      pipeline_EXMEM_stage_N45, pipeline_EXMEM_stage_N44, 
      pipeline_EXMEM_stage_N43, pipeline_EXMEM_stage_N42, 
      pipeline_EXMEM_stage_N41, pipeline_EXMEM_stage_N40, 
      pipeline_EXMEM_stage_N39, pipeline_EXMEM_stage_N38, 
      pipeline_EXMEM_stage_N37, pipeline_EXMEM_stage_N36, 
      pipeline_EXMEM_stage_N35, pipeline_EXMEM_stage_N34, 
      pipeline_EXMEM_stage_N33, pipeline_EXMEM_stage_N32, 
      pipeline_EXMEM_stage_N31, pipeline_EXMEM_stage_N30, 
      pipeline_EXMEM_stage_N29, pipeline_EXMEM_stage_N28, 
      pipeline_EXMEM_stage_N27, pipeline_EXMEM_stage_N26, 
      pipeline_EXMEM_stage_N25, pipeline_EXMEM_stage_N24, 
      pipeline_EXMEM_stage_N23, pipeline_EXMEM_stage_N22, 
      pipeline_EXMEM_stage_N21, pipeline_EXMEM_stage_N20, 
      pipeline_EXMEM_stage_N19, pipeline_EXMEM_stage_N18, 
      pipeline_EXMEM_stage_N17, pipeline_EXMEM_stage_N16, 
      pipeline_EXMEM_stage_N15, pipeline_EXMEM_stage_N14, 
      pipeline_EXMEM_stage_N13, pipeline_EXMEM_stage_N12, 
      pipeline_EXMEM_stage_N11, pipeline_EXMEM_stage_N10, 
      pipeline_EXMEM_stage_N9, pipeline_EXMEM_stage_N8, pipeline_EXMEM_stage_N7
      , pipeline_EXMEM_stage_N6, pipeline_EXMEM_stage_N5, 
      pipeline_EXMEM_stage_N4, pipeline_EXMEM_stage_N3, 
      pipeline_MEMWB_Stage_N47, pipeline_MEMWB_Stage_N46, 
      pipeline_MEMWB_Stage_N45, pipeline_MEMWB_Stage_N44, 
      pipeline_MEMWB_Stage_N43, pipeline_MEMWB_Stage_N42, 
      pipeline_MEMWB_Stage_N41, pipeline_MEMWB_Stage_N40, 
      pipeline_MEMWB_Stage_N39, pipeline_MEMWB_Stage_N38, 
      pipeline_MEMWB_Stage_N37, pipeline_MEMWB_Stage_N36, 
      pipeline_MEMWB_Stage_N35, pipeline_MEMWB_Stage_N34, 
      pipeline_MEMWB_Stage_N33, pipeline_MEMWB_Stage_N32, 
      pipeline_MEMWB_Stage_N31, pipeline_MEMWB_Stage_N30, 
      pipeline_MEMWB_Stage_N29, pipeline_MEMWB_Stage_N28, 
      pipeline_MEMWB_Stage_N27, pipeline_MEMWB_Stage_N26, 
      pipeline_MEMWB_Stage_N25, pipeline_MEMWB_Stage_N24, 
      pipeline_MEMWB_Stage_N23, pipeline_MEMWB_Stage_N22, 
      pipeline_MEMWB_Stage_N21, pipeline_MEMWB_Stage_N20, 
      pipeline_MEMWB_Stage_N19, pipeline_MEMWB_Stage_N18, 
      pipeline_MEMWB_Stage_N17, pipeline_MEMWB_Stage_N16, 
      pipeline_MEMWB_Stage_N15, pipeline_MEMWB_Stage_N14, 
      pipeline_MEMWB_Stage_N13, pipeline_MEMWB_Stage_N12, 
      pipeline_MEMWB_Stage_N11, pipeline_MEMWB_Stage_N10, 
      pipeline_cu_hazard_N40, pipeline_cu_hazard_N39, pipeline_cu_pipeline_N113
      , pipeline_cu_pipeline_N112, pipeline_cu_pipeline_N110, 
      pipeline_cu_pipeline_N109, pipeline_cu_pipeline_N108, 
      pipeline_cu_pipeline_N107, pipeline_cu_pipeline_N106, 
      pipeline_cu_pipeline_N105, pipeline_cu_pipeline_N104, 
      pipeline_cu_pipeline_N103, pipeline_cu_pipeline_N102, 
      pipeline_cu_pipeline_N101, pipeline_cu_pipeline_N89, 
      pipeline_cu_pipeline_N88, DataMem_N2349, DataMem_N2346, DataMem_N2343, 
      DataMem_N2340, DataMem_N2337, DataMem_N2334, DataMem_N2331, DataMem_N2328
      , DataMem_N2325, DataMem_N2322, DataMem_N2319, DataMem_N2316, 
      DataMem_N2313, DataMem_N2310, DataMem_N2307, DataMem_N2304, DataMem_N2301
      , DataMem_N2298, DataMem_N2295, DataMem_N2292, DataMem_N2289, 
      DataMem_N2286, DataMem_N2283, DataMem_N2280, DataMem_N2277, DataMem_N2274
      , DataMem_N2271, DataMem_N2268, DataMem_N2265, DataMem_N2262, 
      DataMem_N2259, DataMem_N2256, DataMem_N2254, DataMem_N2251, DataMem_N2248
      , DataMem_N2245, DataMem_N2242, DataMem_N2239, DataMem_N2236, 
      DataMem_N2233, DataMem_N2230, DataMem_N2227, DataMem_N2224, DataMem_N2221
      , DataMem_N2218, DataMem_N2215, DataMem_N2212, DataMem_N2209, 
      DataMem_N2206, DataMem_N2203, DataMem_N2200, DataMem_N2197, DataMem_N2194
      , DataMem_N2191, DataMem_N2188, DataMem_N2185, DataMem_N2182, 
      DataMem_N2179, DataMem_N2176, DataMem_N2173, DataMem_N2170, DataMem_N2167
      , DataMem_N2164, DataMem_N2161, DataMem_N2159, DataMem_N2157, 
      DataMem_N2155, DataMem_N2153, DataMem_N2151, DataMem_N2149, DataMem_N2147
      , DataMem_N2145, DataMem_N2143, DataMem_N2141, DataMem_N2139, 
      DataMem_N2137, DataMem_N2135, DataMem_N2133, DataMem_N2131, DataMem_N2129
      , DataMem_N2127, DataMem_N2125, DataMem_N2123, DataMem_N2121, 
      DataMem_N2119, DataMem_N2117, DataMem_N2115, DataMem_N2113, DataMem_N2111
      , DataMem_N2109, DataMem_N2107, DataMem_N2105, DataMem_N2103, 
      DataMem_N2101, DataMem_N2099, DataMem_N2097, DataMem_N2095, DataMem_N2093
      , DataMem_N2091, DataMem_N2089, DataMem_N2087, DataMem_N2085, 
      DataMem_N2083, DataMem_N2081, DataMem_N2079, DataMem_N2077, DataMem_N2075
      , DataMem_N2073, DataMem_N2071, DataMem_N2069, DataMem_N2067, 
      DataMem_N2065, DataMem_N2063, DataMem_N2061, DataMem_N2059, DataMem_N2057
      , DataMem_N2055, DataMem_N2053, DataMem_N2051, DataMem_N2049, 
      DataMem_N2047, DataMem_N2045, DataMem_N2043, DataMem_N2041, DataMem_N2039
      , DataMem_N2037, DataMem_N2035, DataMem_N2033, DataMem_N2031, 
      DataMem_N2029, DataMem_N2027, DataMem_N2025, DataMem_N2023, DataMem_N2021
      , DataMem_N2019, DataMem_N2017, DataMem_N2015, DataMem_N2013, 
      DataMem_N2011, DataMem_N2009, DataMem_N2007, DataMem_N2005, DataMem_N2003
      , DataMem_N2001, DataMem_N1999, DataMem_N1997, DataMem_N1995, 
      DataMem_N1993, DataMem_N1991, DataMem_N1989, DataMem_N1987, DataMem_N1985
      , DataMem_N1983, DataMem_N1981, DataMem_N1979, DataMem_N1977, 
      DataMem_N1975, DataMem_N1973, DataMem_N1971, DataMem_N1969, DataMem_N1967
      , DataMem_N1965, DataMem_N1963, DataMem_N1961, DataMem_N1959, 
      DataMem_N1957, DataMem_N1955, DataMem_N1953, DataMem_N1951, DataMem_N1949
      , DataMem_N1947, DataMem_N1945, DataMem_N1943, DataMem_N1941, 
      DataMem_N1939, DataMem_N1937, DataMem_N1935, DataMem_N1933, DataMem_N1931
      , DataMem_N1929, DataMem_N1927, DataMem_N1925, DataMem_N1923, 
      DataMem_N1921, DataMem_N1919, DataMem_N1917, DataMem_N1915, DataMem_N1913
      , DataMem_N1911, DataMem_N1909, DataMem_N1907, DataMem_N1905, 
      DataMem_N1903, DataMem_N1901, DataMem_N1899, DataMem_N1897, DataMem_N1895
      , DataMem_N1893, DataMem_N1891, DataMem_N1889, DataMem_N1887, 
      DataMem_N1885, DataMem_N1883, DataMem_N1881, DataMem_N1879, DataMem_N1877
      , DataMem_N1875, DataMem_N1873, DataMem_N1871, DataMem_N1869, 
      DataMem_N1867, DataMem_N1865, DataMem_N1863, DataMem_N1861, DataMem_N1859
      , DataMem_N1857, DataMem_N1855, DataMem_N1853, DataMem_N1851, 
      DataMem_N1849, DataMem_N1847, DataMem_N1845, DataMem_N1843, DataMem_N1841
      , DataMem_N1839, DataMem_N1837, DataMem_N1835, DataMem_N1833, 
      DataMem_N1831, DataMem_N1829, DataMem_N1827, DataMem_N1825, DataMem_N1823
      , DataMem_N1821, DataMem_N1819, DataMem_N1817, DataMem_N1815, 
      DataMem_N1813, DataMem_N1811, DataMem_N1809, DataMem_N1807, DataMem_N1805
      , DataMem_N1803, DataMem_N1801, DataMem_N1799, DataMem_N1797, 
      DataMem_N1795, DataMem_N1793, DataMem_N1791, DataMem_N1789, DataMem_N1787
      , DataMem_N1785, DataMem_N1783, DataMem_N1781, DataMem_N1779, 
      DataMem_N1777, DataMem_N1775, DataMem_N1773, DataMem_N1771, DataMem_N1769
      , DataMem_N1767, DataMem_N1765, DataMem_N1763, DataMem_N1761, 
      DataMem_N1759, DataMem_N1757, DataMem_N1755, DataMem_N1753, DataMem_N1751
      , DataMem_N1749, DataMem_N1747, DataMem_N1745, DataMem_N1743, 
      DataMem_N1741, DataMem_N1739, DataMem_N1737, DataMem_N1735, DataMem_N1733
      , DataMem_N1731, DataMem_N1729, DataMem_N1727, DataMem_N1725, 
      DataMem_N1723, DataMem_N1721, DataMem_N1719, DataMem_N1717, DataMem_N1715
      , DataMem_N1713, DataMem_N1711, DataMem_N1709, DataMem_N1707, 
      DataMem_N1705, DataMem_N1703, DataMem_N1701, DataMem_N1699, DataMem_N1697
      , DataMem_N1695, DataMem_N1693, DataMem_N1691, DataMem_N1689, 
      DataMem_N1687, DataMem_N1685, DataMem_N1683, DataMem_N1681, DataMem_N1679
      , DataMem_N1677, DataMem_N1675, DataMem_N1673, DataMem_N1671, 
      DataMem_N1669, DataMem_N1667, DataMem_N1665, DataMem_N1663, DataMem_N1661
      , DataMem_N1659, DataMem_N1657, DataMem_N1655, DataMem_N1653, 
      DataMem_N1651, DataMem_N1649, DataMem_Mem_0_0_port, DataMem_Mem_0_1_port,
      DataMem_Mem_0_2_port, DataMem_Mem_0_3_port, DataMem_Mem_0_4_port, 
      DataMem_Mem_0_5_port, DataMem_Mem_0_6_port, DataMem_Mem_0_7_port, 
      DataMem_Mem_0_8_port, DataMem_Mem_0_9_port, DataMem_Mem_0_10_port, 
      DataMem_Mem_0_11_port, DataMem_Mem_0_12_port, DataMem_Mem_0_13_port, 
      DataMem_Mem_0_14_port, DataMem_Mem_0_15_port, DataMem_Mem_0_16_port, 
      DataMem_Mem_0_17_port, DataMem_Mem_0_18_port, DataMem_Mem_0_19_port, 
      DataMem_Mem_0_20_port, DataMem_Mem_0_21_port, DataMem_Mem_0_22_port, 
      DataMem_Mem_0_23_port, DataMem_Mem_0_24_port, DataMem_Mem_0_25_port, 
      DataMem_Mem_0_26_port, DataMem_Mem_0_27_port, DataMem_Mem_0_28_port, 
      DataMem_Mem_0_29_port, DataMem_Mem_0_30_port, DataMem_Mem_0_31_port, 
      DataMem_Mem_1_0_port, DataMem_Mem_1_1_port, DataMem_Mem_1_2_port, 
      DataMem_Mem_1_3_port, DataMem_Mem_1_4_port, DataMem_Mem_1_5_port, 
      DataMem_Mem_1_6_port, DataMem_Mem_1_7_port, DataMem_Mem_1_8_port, 
      DataMem_Mem_1_9_port, DataMem_Mem_1_10_port, DataMem_Mem_1_11_port, 
      DataMem_Mem_1_12_port, DataMem_Mem_1_13_port, DataMem_Mem_1_14_port, 
      DataMem_Mem_1_15_port, DataMem_Mem_1_16_port, DataMem_Mem_1_17_port, 
      DataMem_Mem_1_18_port, DataMem_Mem_1_19_port, DataMem_Mem_1_20_port, 
      DataMem_Mem_1_21_port, DataMem_Mem_1_22_port, DataMem_Mem_1_23_port, 
      DataMem_Mem_1_24_port, DataMem_Mem_1_25_port, DataMem_Mem_1_26_port, 
      DataMem_Mem_1_27_port, DataMem_Mem_1_28_port, DataMem_Mem_1_29_port, 
      DataMem_Mem_1_30_port, DataMem_Mem_1_31_port, DataMem_Mem_2_0_port, 
      DataMem_Mem_2_1_port, DataMem_Mem_2_2_port, DataMem_Mem_2_3_port, 
      DataMem_Mem_2_4_port, DataMem_Mem_2_5_port, DataMem_Mem_2_6_port, 
      DataMem_Mem_2_7_port, DataMem_Mem_2_8_port, DataMem_Mem_2_9_port, 
      DataMem_Mem_2_10_port, DataMem_Mem_2_11_port, DataMem_Mem_2_12_port, 
      DataMem_Mem_2_13_port, DataMem_Mem_2_14_port, DataMem_Mem_2_15_port, 
      DataMem_Mem_2_16_port, DataMem_Mem_2_17_port, DataMem_Mem_2_18_port, 
      DataMem_Mem_2_19_port, DataMem_Mem_2_20_port, DataMem_Mem_2_21_port, 
      DataMem_Mem_2_22_port, DataMem_Mem_2_23_port, DataMem_Mem_2_24_port, 
      DataMem_Mem_2_25_port, DataMem_Mem_2_26_port, DataMem_Mem_2_27_port, 
      DataMem_Mem_2_28_port, DataMem_Mem_2_29_port, DataMem_Mem_2_30_port, 
      DataMem_Mem_2_31_port, DataMem_Mem_3_0_port, DataMem_Mem_3_1_port, 
      DataMem_Mem_3_2_port, DataMem_Mem_3_3_port, DataMem_Mem_3_4_port, 
      DataMem_Mem_3_5_port, DataMem_Mem_3_6_port, DataMem_Mem_3_7_port, 
      DataMem_Mem_3_8_port, DataMem_Mem_3_9_port, DataMem_Mem_3_10_port, 
      DataMem_Mem_3_11_port, DataMem_Mem_3_12_port, DataMem_Mem_3_13_port, 
      DataMem_Mem_3_14_port, DataMem_Mem_3_15_port, DataMem_Mem_3_16_port, 
      DataMem_Mem_3_17_port, DataMem_Mem_3_18_port, DataMem_Mem_3_19_port, 
      DataMem_Mem_3_20_port, DataMem_Mem_3_21_port, DataMem_Mem_3_22_port, 
      DataMem_Mem_3_23_port, DataMem_Mem_3_24_port, DataMem_Mem_3_25_port, 
      DataMem_Mem_3_26_port, DataMem_Mem_3_27_port, DataMem_Mem_3_28_port, 
      DataMem_Mem_3_29_port, DataMem_Mem_3_30_port, DataMem_Mem_3_31_port, 
      DataMem_Mem_4_0_port, DataMem_Mem_4_1_port, DataMem_Mem_4_2_port, 
      DataMem_Mem_4_3_port, DataMem_Mem_4_4_port, DataMem_Mem_4_5_port, 
      DataMem_Mem_4_6_port, DataMem_Mem_4_7_port, DataMem_Mem_4_8_port, 
      DataMem_Mem_4_9_port, DataMem_Mem_4_10_port, DataMem_Mem_4_11_port, 
      DataMem_Mem_4_12_port, DataMem_Mem_4_13_port, DataMem_Mem_4_14_port, 
      DataMem_Mem_4_15_port, DataMem_Mem_4_16_port, DataMem_Mem_4_17_port, 
      DataMem_Mem_4_18_port, DataMem_Mem_4_19_port, DataMem_Mem_4_20_port, 
      DataMem_Mem_4_21_port, DataMem_Mem_4_22_port, DataMem_Mem_4_23_port, 
      DataMem_Mem_4_24_port, DataMem_Mem_4_25_port, DataMem_Mem_4_26_port, 
      DataMem_Mem_4_27_port, DataMem_Mem_4_28_port, DataMem_Mem_4_29_port, 
      DataMem_Mem_4_30_port, DataMem_Mem_4_31_port, DataMem_Mem_5_0_port, 
      DataMem_Mem_5_1_port, DataMem_Mem_5_2_port, DataMem_Mem_5_3_port, 
      DataMem_Mem_5_4_port, DataMem_Mem_5_5_port, DataMem_Mem_5_6_port, 
      DataMem_Mem_5_7_port, DataMem_Mem_5_8_port, DataMem_Mem_5_9_port, 
      DataMem_Mem_5_10_port, DataMem_Mem_5_11_port, DataMem_Mem_5_12_port, 
      DataMem_Mem_5_13_port, DataMem_Mem_5_14_port, DataMem_Mem_5_15_port, 
      DataMem_Mem_5_16_port, DataMem_Mem_5_17_port, DataMem_Mem_5_18_port, 
      DataMem_Mem_5_19_port, DataMem_Mem_5_20_port, DataMem_Mem_5_21_port, 
      DataMem_Mem_5_22_port, DataMem_Mem_5_23_port, DataMem_Mem_5_24_port, 
      DataMem_Mem_5_25_port, DataMem_Mem_5_26_port, DataMem_Mem_5_27_port, 
      DataMem_Mem_5_28_port, DataMem_Mem_5_29_port, DataMem_Mem_5_30_port, 
      DataMem_Mem_5_31_port, DataMem_Mem_6_0_port, DataMem_Mem_6_1_port, 
      DataMem_Mem_6_2_port, DataMem_Mem_6_3_port, DataMem_Mem_6_4_port, 
      DataMem_Mem_6_5_port, DataMem_Mem_6_6_port, DataMem_Mem_6_7_port, 
      DataMem_Mem_6_8_port, DataMem_Mem_6_9_port, DataMem_Mem_6_10_port, 
      DataMem_Mem_6_11_port, DataMem_Mem_6_12_port, DataMem_Mem_6_13_port, 
      DataMem_Mem_6_14_port, DataMem_Mem_6_15_port, DataMem_Mem_6_16_port, 
      DataMem_Mem_6_17_port, DataMem_Mem_6_18_port, DataMem_Mem_6_19_port, 
      DataMem_Mem_6_20_port, DataMem_Mem_6_21_port, DataMem_Mem_6_22_port, 
      DataMem_Mem_6_23_port, DataMem_Mem_6_24_port, DataMem_Mem_6_25_port, 
      DataMem_Mem_6_26_port, DataMem_Mem_6_27_port, DataMem_Mem_6_28_port, 
      DataMem_Mem_6_29_port, DataMem_Mem_6_30_port, DataMem_Mem_6_31_port, 
      DataMem_Mem_7_0_port, DataMem_Mem_7_1_port, DataMem_Mem_7_2_port, 
      DataMem_Mem_7_3_port, DataMem_Mem_7_4_port, DataMem_Mem_7_5_port, 
      DataMem_Mem_7_6_port, DataMem_Mem_7_7_port, DataMem_Mem_7_8_port, 
      DataMem_Mem_7_9_port, DataMem_Mem_7_10_port, DataMem_Mem_7_11_port, 
      DataMem_Mem_7_12_port, DataMem_Mem_7_13_port, DataMem_Mem_7_14_port, 
      DataMem_Mem_7_15_port, DataMem_Mem_7_16_port, DataMem_Mem_7_17_port, 
      DataMem_Mem_7_18_port, DataMem_Mem_7_19_port, DataMem_Mem_7_20_port, 
      DataMem_Mem_7_21_port, DataMem_Mem_7_22_port, DataMem_Mem_7_23_port, 
      DataMem_Mem_7_24_port, DataMem_Mem_7_25_port, DataMem_Mem_7_26_port, 
      DataMem_Mem_7_27_port, DataMem_Mem_7_28_port, DataMem_Mem_7_29_port, 
      DataMem_Mem_7_30_port, DataMem_Mem_7_31_port, DataMem_N31, DataMem_N30, 
      DataMem_N29, DataMem_N28, DataMem_N27, DataMem_N26, DataMem_N25, 
      DataMem_N24, DataMem_N23, DataMem_N22, DataMem_N21, DataMem_N20, 
      DataMem_N19, DataMem_N18, DataMem_N17, DataMem_N16, DataMem_N15, 
      DataMem_N14, DataMem_N13, DataMem_N12, DataMem_N11, DataMem_N10, 
      DataMem_N9, DataMem_N8, DataMem_N7, DataMem_N6, DataMem_N5, DataMem_N4, 
      DataMem_N3, DataMem_N2, DataMem_N1, DataMem_N0, n415, n3855, n3856, n3857
      , n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, 
      n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, 
      n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, 
      n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, 
      n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, 
      n3908, n3909, n3910, n3911, n3912, n3923, n3924, n3925, n3926, n3927, 
      n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, 
      n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, 
      n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, 
      n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, 
      n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, 
      n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, 
      n3988, n3989, n3990, n3991, n3992, n4376, n7648, n7649, n7650, n7651, 
      n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, 
      n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, 
      n7672, n7673, n7674, n7675, n7676, n7709, n7710, n7711, net175543, n12625
      , n12649, n12766, n13055, n13058, n13061, n13064, n13067, n13070, n13073,
      n13076, n13079, n13082, n13085, n13088, n13091, n13094, n13097, n13100, 
      n13103, n13106, n13109, n13112, n13115, n13118, n13121, n13124, n13127, 
      n13130, n13133, n13136, n13139, n13142, n13145, n13148, n13151, n13154, 
      n13157, n13160, n13163, n13166, n13169, n13172, n13175, n13178, n13181, 
      n13184, n13187, n13190, n13193, n13196, n13199, n13202, n13205, n13208, 
      n13211, n13214, n13217, n13220, n13223, n13226, n13229, n13232, n13235, 
      n13238, n13241, n13244, n13247, n13250, n13253, n13256, n13259, n13262, 
      n13265, n13268, n13782, n13783, n13784, n13785, n13786, n13787, n13788, 
      n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797, 
      n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806, 
      n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815, 
      n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824, 
      n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833, 
      n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842, 
      n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851, 
      n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860, 
      n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869, 
      n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878, 
      n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13925, 
      n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934, 
      n13936, n13937, n13938, n13939, n13940, n13942, n13944, n13945, n13946, 
      n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955, 
      n13956, n13957, n13958, n13959, n13960, n13962, n13963, n13964, n13965, 
      n13966, n13967, n13969, n13979, n13980, n13981, n13982, n13983, n13984, 
      n13985, n13986, n13987, n13988, n13989, n13990, n13992, n13993, n13994, 
      n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003, 
      n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012, 
      n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021, 
      n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030, 
      n14031, n14032, n14033, n14034, n14035, n14040, n14041, n14042, n14043, 
      n14044, n14045, n14046, n14047, n14048, n14049, n14051, n14053, n14058, 
      n14059, n14061, n14064, n14065, n14066, n14067, n14068, n14069, n14070, 
      n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14082, 
      n14083, n14084, n14086, n14087, n14088, n14089, n14090, n14091, n14092, 
      n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101, 
      n14102, n14103, n14104, n14105, n14113, n14116, n14117, n14119, n14120, 
      n14121, n14122, n14123, n14125, n14126, n14127, n14129, n14133, n14134, 
      n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143, 
      n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152, 
      n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161, 
      n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170, 
      n14172, n14173, n14174, n14176, n14177, n14178, n14179, n14180, n14181, 
      n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14200, 
      n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14210, 
      n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220, 
      n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229, 
      n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238, 
      n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247, 
      n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256, 
      n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265, 
      n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274, 
      n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283, 
      n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292, 
      n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301, 
      n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310, 
      n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319, 
      n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328, 
      n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337, 
      n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346, 
      n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355, 
      n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364, 
      n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373, 
      n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382, 
      n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391, 
      n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400, 
      n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409, 
      n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418, 
      n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427, 
      n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436, 
      n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445, 
      n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454, 
      n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463, 
      n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472, 
      n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481, 
      n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490, 
      n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499, 
      n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508, 
      n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517, 
      n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526, 
      n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535, 
      n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544, 
      n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553, 
      n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562, 
      n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571, 
      n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580, 
      n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589, 
      n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598, 
      n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607, 
      n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616, 
      n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625, 
      n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634, 
      n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643, 
      n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652, 
      n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661, 
      n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670, 
      n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679, 
      n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688, 
      n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697, 
      n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706, 
      n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715, 
      n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724, 
      n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733, 
      n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742, 
      n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751, 
      n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760, 
      n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769, 
      n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778, 
      n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787, 
      n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796, 
      n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805, 
      n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814, 
      n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823, 
      n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832, 
      n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841, 
      n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850, 
      n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859, 
      n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868, 
      n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877, 
      n14878, n14879, n14880, n14881, n14882, n14883, n14885, n14887, n14889, 
      n14891, n14893, n14895, n14897, n14899, n14901, n14903, n14905, n14907, 
      n14909, n14911, n14913, n14915, n14917, n14919, n14921, n14923, n14925, 
      n14927, n14929, n14931, n14933, n14935, n14937, n14939, n14941, n14943, 
      n14945, n14947, n14948, n14949, n14950, n14951, n14952, n14954, n14955, 
      n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964, 
      n14965, n14966, n14967, n14968, n14970, n14971, n14972, n14974, n14975, 
      n14976, n14977, n14978, n14979, n14981, n14982, n14988, n14993, n14995, 
      n15001, n15007, n15009, n15010, n15011, n15013, n15014, n15015, n15017, 
      n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15029, 
      n15030, n15032, n15033, n15034, n15035, n15037, n15039, n15040, n15041, 
      n15042, n15043, n15045, n15046, n15047, n15048, n15049, n15050, n15051, 
      n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15062, n15064, 
      n15066, n15068, n15070, n15072, n15074, n15076, n15078, n15080, n15082, 
      n15084, n15086, n15088, n15090, n15092, n15094, n15096, n15098, n15100, 
      n15102, n15104, n15106, n15108, n15110, n15112, n15114, n15116, n15118, 
      n15120, n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129, 
      n15130, n15131, n15133, n15134, n15137, n15138, n15142, n15145, n15146, 
      n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155, 
      n15156, n15157, n15159, n15160, n15161, n15162, n15163, n15164, n15165, 
      n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174, 
      n15175, n15176, n15180, n15181, n15182, n15183, n15184, n15185, n15186, 
      n15187, n15188, n15189, n15191, n15192, n15193, n15194, n15195, n15196, 
      n15197, n15198, n15199, n15201, n15202, n15204, n15205, n15206, n15207, 
      n15208, n15209, n15210, n15211, n15212, n15213, n15215, n15216, n15217, 
      n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226, 
      n15227, n15228, n15229, n15230, n15231, n15233, n15234, n15235, n15236, 
      n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15245, n15246, 
      n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255, 
      n15256, n15257, n15258, n15260, n15261, n15262, n15263, n15264, n15265, 
      n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274, 
      n15275, n15276, n15278, n15279, n15280, n15281, n15282, n15283, n15284, 
      n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15294, 
      n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303, 
      n15304, n15305, n15306, n15307, n15308, n15309, n15311, n15312, n15313, 
      n15314, n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323, 
      n15324, n15325, n15326, n15327, n15328, n15330, n15331, n15332, n15333, 
      n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342, 
      n15343, n15345, n15346, n15348, n15352, n15353, n15354, n15355, n15356, 
      n15357, n15358, n15359, n15360, n15362, n15363, n15366, n15367, n15368, 
      n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377, 
      n15378, n15379, n15381, n15382, n15383, n15384, n15385, n15386, n15387, 
      n15388, n15389, n15390, n15391, n15392, n15393, n15395, n15396, n15397, 
      n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406, 
      n15407, n15408, n15410, n15411, n15412, n15413, n15414, n15415, n15416, 
      n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425, 
      n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434, 
      n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15444, 
      n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453, 
      n15454, n15455, n15456, n15458, n15459, n15460, n15461, n15462, n15463, 
      n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15473, 
      n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15482, n15483, 
      n15484, n15485, n15486, n15487, n15488, n15489, n15491, n15492, n15493, 
      n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502, 
      n15503, n15504, n15505, n15507, n15508, n15509, n15510, n15511, n15512, 
      n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15521, n15522, 
      n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531, 
      n15532, n15533, n15534, n15535, n15537, n15538, n15539, n15540, n15541, 
      n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550, 
      n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560, 
      n15561, n15562, n15563, n15564, n15566, n15567, n15568, n15569, n15570, 
      n15571, n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15581, 
      n15582, n15583, n15584, n15586, n15588, n15590, n15591, n15592, n15593, 
      n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602, 
      n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611, 
      n15612, n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628, 
      n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637, 
      n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646, 
      n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15686, n15687, 
      n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696, 
      n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705, 
      n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714, 
      n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723, 
      n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732, 
      n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741, 
      n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750, 
      n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759, 
      n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768, 
      n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777, 
      n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786, 
      n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795, 
      n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804, 
      n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813, 
      n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822, 
      n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831, 
      n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840, 
      n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849, 
      n15866, n15867, n15868, n15869, n15886, n15887, n15888, n15889, n15890, 
      n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899, 
      n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909, 
      n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917, n15918, 
      n15919, n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927, 
      n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936, 
      n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945, 
      n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954, 
      n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963, 
      n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972, 
      n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981, 
      n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989, n15990, 
      n15991, n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999, 
      n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008, 
      n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017, 
      n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026, 
      n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035, 
      n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043, n16044, 
      n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053, 
      n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061, n16062, 
      n16063, n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071, 
      n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080, 
      n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089, 
      n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098, 
      n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107, 
      n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115, n16116, 
      n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125, 
      n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133, n16134, 
      n16135, n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143, 
      n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152, 
      n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161, 
      n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170, 
      n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179, 
      n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187, n16188, 
      n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197, 
      n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205, n16206, 
      n16207, n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215, 
      n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224, 
      n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233, 
      n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242, 
      n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251, 
      n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259, n16260, 
      n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269, 
      n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277, n16278, 
      n16279, n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287, 
      n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296, 
      n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305, 
      n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314, 
      n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323, 
      n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332, 
      n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341, 
      n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349, n16350, 
      n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359, 
      n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368, 
      n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377, 
      n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386, 
      n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395, 
      n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404, 
      n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413, 
      n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421, n16422, 
      n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431, 
      n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440, 
      n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449, 
      n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458, 
      n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467, 
      n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476, 
      n16477, n16478, n16479, n16480, n16481, n16482, n16483, n16484, n16485, 
      n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16493, n16494, 
      n16495, n16496, n16497, n16498, n16499, n16500, n16501, n16502, n16503, 
      n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512, 
      n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521, 
      n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530, 
      n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539, 
      n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548, 
      n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556, n16557, 
      n16558, n16559, n16560, n16561, n16562, n16563, n16565, n16568, n16571, 
      n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580, 
      n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588, n16589, 
      n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597, n16598, 
      n16599, n16603, n16605, n16606, n16607, n16608, n16609, n16611, n16612, 
      n16614, n16615, n16616, n16617, n16618, n16619, n16620, n16624, n16626, 
      n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637, 
      n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645, n16646, 
      n16647, n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655, 
      n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664, 
      n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16676, n16677, 
      n16678, n16679, n16680, n16681, n16683, n16684, n16685, n16686, n16687, 
      n16689, n16690, n16691, n16693, n16696, n16699, n16701, n16704, n16710, 
      n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719, 
      n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728, 
      n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737, 
      n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746, 
      n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755, 
      n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764, 
      n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772, n16773, 
      n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16784, n16785, 
      n16786, n16789, n16790, n16791, n16792, n16793, n16795, n16796, n16806, 
      n16807, n16808, n16809, n16811, n16812, n16813, n16814, n16815, n16816, 
      n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825, 
      n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834, 
      n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843, 
      n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851, n16852, 
      n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860, n16861, 
      n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869, n16870, 
      n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879, 
      n16880, n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888, 
      n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897, 
      n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906, 
      n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915, 
      n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923, n16924, 
      n16925, n16926, n16927, n16928, n16929, n16930, n16931, n16932, n16933, 
      n16934, n16935, n16936, n16937, n16938, n16939, n16940, n16941, n16942, 
      n16943, n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951, 
      n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960, 
      n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969, 
      n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978, 
      n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987, 
      n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995, n16996, 
      n16997, n16998, n16999, n17000, n17001, n17002, n17003, n17004, n17005, 
      n17006, n17007, n17008, n17009, n17010, n17011, n17012, n17013, n17014, 
      n17015, n17016, n16613, n16682, n16688, n16805, n15000, n16783, n16782, 
      n15005, pipeline_stageF_PC_plus4_add_26_n1, 
      pipeline_stageF_PC_plus4_add_26_carry_4_port, 
      pipeline_stageF_PC_plus4_add_26_carry_5_port, 
      pipeline_stageF_PC_plus4_add_26_carry_6_port, 
      pipeline_stageF_PC_plus4_add_26_carry_7_port, 
      pipeline_stageF_PC_plus4_add_26_carry_8_port, 
      pipeline_stageF_PC_plus4_add_26_carry_9_port, 
      pipeline_stageF_PC_plus4_add_26_carry_10_port, 
      pipeline_stageF_PC_plus4_add_26_carry_11_port, 
      pipeline_stageF_PC_plus4_add_26_carry_12_port, 
      pipeline_stageF_PC_plus4_add_26_carry_13_port, 
      pipeline_stageF_PC_plus4_add_26_carry_14_port, 
      pipeline_stageF_PC_plus4_add_26_carry_15_port, 
      pipeline_stageF_PC_plus4_add_26_carry_16_port, 
      pipeline_stageF_PC_plus4_add_26_carry_17_port, 
      pipeline_stageF_PC_plus4_add_26_carry_18_port, 
      pipeline_stageF_PC_plus4_add_26_carry_19_port, 
      pipeline_stageF_PC_plus4_add_26_carry_20_port, 
      pipeline_stageF_PC_plus4_add_26_carry_21_port, 
      pipeline_stageF_PC_plus4_add_26_carry_22_port, 
      pipeline_stageF_PC_plus4_add_26_carry_23_port, 
      pipeline_stageF_PC_plus4_add_26_carry_24_port, 
      pipeline_stageF_PC_plus4_add_26_carry_25_port, 
      pipeline_stageF_PC_plus4_add_26_carry_26_port, 
      pipeline_stageF_PC_plus4_add_26_carry_27_port, 
      pipeline_stageF_PC_plus4_add_26_carry_28_port, 
      pipeline_stageF_PC_plus4_add_26_carry_29_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n170, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n169, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n167, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n166, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n165, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n164, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n163, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n162, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n161, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n160, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n158, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n157, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n156, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n155, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n154, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n153, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n152, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n151, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n150, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n149, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n148, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n145, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n144, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n143, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n140, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n139, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n136, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n135, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n134, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n133, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n132, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n127, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n124, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n121, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n118, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n117, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n116, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n115, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n114, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n113, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n112, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n111, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n110, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n109, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n108, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n107, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n106, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n105, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n103, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n102, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n101, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n100, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n99, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n98, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n94, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n93, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n92, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n91, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n90, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n89, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n88, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n87, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n86, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n85, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n84, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n83, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n82, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n81, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n80, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n79, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n78, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n77, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n76, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n75, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n74, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n73, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n72, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n71, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n70, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n69, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n68, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n67, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n66, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n64, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n63, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n62, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n61, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n60, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n59, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n58, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n56, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n54, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n53, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n52, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n51, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n50, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n48, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n46, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n45, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n44, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n43, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n42, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n41, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n40, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n39, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n38, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n37, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n36, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n35, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n34, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n33, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n32, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n31, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n30, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n29, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n28, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n27, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n26, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n25, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n24, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n23, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n22, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n21, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n20, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n19, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n18, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n17, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n16, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n15, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n14, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n13, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n12, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n11, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n10, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n9, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n8, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n7, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n6, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n5, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n4, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n2, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_n1, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_SH_1_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_SH_3_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C48_A_16_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n172, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n171, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n170, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n169, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n168, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n167, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n165, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n163, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n162, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n161, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n160, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n158, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n156, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n154, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n153, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n152, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n149, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n146, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n144, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n143, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n142, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n140, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n139, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n138, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n136, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n135, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n134, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n133, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n131, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n130, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n129, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n128, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n127, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n126, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n122, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n121, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n120, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n118, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n117, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n116, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n114, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n113, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n112, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n111, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n109, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n108, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n107, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n106, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n104, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n103, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n102, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n101, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n99, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n98, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n97, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n96, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n95, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n94, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n92, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n91, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n90, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n89, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n88, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n87, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n85, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n84, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n83, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n82, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n81, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n80, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n79, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n77, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n76, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n75, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n74, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n73, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n72, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n71, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n70, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n69, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n68, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n67, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n66, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n64, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n63, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n62, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n61, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n60, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n58, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n57, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n56, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n55, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n54, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n53, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n52, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n50, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n49, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n48, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n47, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n46, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n45, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n44, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n42, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n41, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n40, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n39, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n38, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n37, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n36, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n35, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n33, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n32, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n31, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n30, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n29, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n28, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n27, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n26, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n25, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n23, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n21, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n20, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n19, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n18, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n17, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n16, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n15, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n14, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n13, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n12, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n11, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n10, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n9, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n8, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n7, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n6, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n5, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n4, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n3, 
      pipeline_stageE_EXE_ALU_alu_shift_C86_n1, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_0_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_1_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_2_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_3_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_4_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_5_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_6_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_7_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_8_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_9_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_10_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_11_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_12_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_13_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_14_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_15_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_16_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_17_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_18_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_19_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_20_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_21_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_22_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_23_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_24_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_25_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_26_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_27_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_28_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_29_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_30_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_31_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_0_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_1_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_2_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_3_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_4_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_5_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_6_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_7_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_8_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_9_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_10_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_11_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_12_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_13_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_14_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_15_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_16_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_17_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_18_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_19_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_20_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_21_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_22_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_23_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_24_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_25_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_26_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_27_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_28_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_29_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_30_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_31_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_0_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_1_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_2_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_3_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_4_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_5_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_6_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_7_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_8_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_9_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_10_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_11_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_12_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_13_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_14_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_15_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_16_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_17_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_18_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_19_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_20_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_21_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_22_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_23_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_24_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_25_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_26_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_27_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_28_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_29_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_30_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_31_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_0_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_1_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_2_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_3_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_5_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_6_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_7_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_8_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_9_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_10_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_11_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_12_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_13_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_14_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_15_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_16_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_17_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_18_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_19_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_20_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_21_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_22_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_23_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_24_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_25_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_26_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_27_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_28_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_29_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_30_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_31_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_0_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_1_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_2_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_3_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_4_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_5_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_6_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_7_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_8_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_9_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_10_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_11_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_12_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_13_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_14_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_15_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_16_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_17_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_18_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_19_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_20_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_21_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_22_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_23_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_24_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_25_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_26_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_27_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_28_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_29_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_30_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_31_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_0_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_1_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_2_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_3_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_4_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_5_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_6_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_7_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_8_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_9_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_10_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_11_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_12_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_13_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_14_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_15_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_16_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_17_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_18_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_19_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_20_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_21_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_22_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_23_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_24_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_25_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_26_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_27_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_28_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_29_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_30_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_31_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_0_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_1_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_2_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_3_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_4_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_5_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_6_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_7_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_8_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_9_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_10_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_11_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_12_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_13_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_14_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_15_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_16_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_17_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_18_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_19_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_20_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_21_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_22_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_23_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_24_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_25_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_26_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_27_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_28_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_29_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_30_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_31_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_0_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_1_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_2_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_3_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_4_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_5_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_6_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_7_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_8_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_9_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_10_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_11_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_12_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_13_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_14_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_15_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_16_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_17_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_18_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_19_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_20_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_21_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_22_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_23_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_24_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_25_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_26_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_27_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_28_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_29_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_30_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_31_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n167, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n161, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n160, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n159, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n158, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n157, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n156, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n155, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n153, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n151, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n148, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n147, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n146, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n145, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n144, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n143, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n142, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n141, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n139, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n138, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n137, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n132, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n131, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n128, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n127, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n126, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n125, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n124, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n123, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n122, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n121, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n120, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n117, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n114, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n108, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n105, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n104, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n103, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n102, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n101, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n100, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n99, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n98, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n97, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n96, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n95, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n94, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n93, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n92, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n91, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n90, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n89, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n88, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n87, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n83, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n82, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n81, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n80, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n79, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n78, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n77, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n76, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n75, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n74, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n73, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n72, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n71, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n70, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n69, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n68, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n67, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n66, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n65, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n63, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n62, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n61, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n60, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n59, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n58, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n57, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n55, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n53, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n51, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n50, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n49, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n48, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n46, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n44, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n43, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n42, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n41, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n40, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n39, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n38, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n37, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n36, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n35, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n34, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n33, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n32, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n31, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n30, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n29, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n28, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n27, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n26, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n25, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n24, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n23, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n22, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n21, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n20, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n19, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n18, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n17, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n16, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n15, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n14, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n13, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n12, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n11, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n10, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n9, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n8, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n7, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n6, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n5, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n4, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n3, 
      pipeline_stageE_EXE_ALU_alu_shift_C50_n2, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_n10, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_n9, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_n8, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_n7, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_n6, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_n5, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_n4, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_n3, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_0_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_1_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_2_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_3_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_4_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_5_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_6_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_7_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_8_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_9_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_10_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_11_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_12_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_13_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_14_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_15_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_16_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_17_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_18_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_19_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_20_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_21_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_22_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_23_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_24_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_25_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_26_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_27_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_28_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_29_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_30_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_31_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_0_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_1_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_2_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_3_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_4_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_5_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_6_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_7_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_8_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_9_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_10_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_11_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_12_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_13_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_14_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_15_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_16_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_17_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_18_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_19_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_20_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_21_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_22_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_23_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_24_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_25_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_26_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_27_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_28_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_29_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_30_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_31_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_0_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_1_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_2_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_3_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_4_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_5_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_6_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_7_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_8_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_9_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_10_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_11_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_12_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_13_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_14_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_15_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_16_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_17_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_18_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_19_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_20_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_21_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_22_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_23_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_24_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_25_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_26_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_27_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_28_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_29_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_30_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_31_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_0_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_1_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_2_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_3_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_4_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_5_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_6_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_7_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_8_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_9_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_10_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_11_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_12_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_13_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_14_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_15_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_16_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_17_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_18_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_19_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_20_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_21_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_22_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_23_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_24_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_25_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_26_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_27_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_28_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_29_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_30_port, 
      pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_31_port, 
      pipeline_stageD_evaluate_jump_target_add_29_n214, 
      pipeline_stageD_evaluate_jump_target_add_29_n213, 
      pipeline_stageD_evaluate_jump_target_add_29_n209, 
      pipeline_stageD_evaluate_jump_target_add_29_n208, 
      pipeline_stageD_evaluate_jump_target_add_29_n207, 
      pipeline_stageD_evaluate_jump_target_add_29_n203, 
      pipeline_stageD_evaluate_jump_target_add_29_n202, 
      pipeline_stageD_evaluate_jump_target_add_29_n201, 
      pipeline_stageD_evaluate_jump_target_add_29_n197, 
      pipeline_stageD_evaluate_jump_target_add_29_n196, 
      pipeline_stageD_evaluate_jump_target_add_29_n195, 
      pipeline_stageD_evaluate_jump_target_add_29_n194, 
      pipeline_stageD_evaluate_jump_target_add_29_n191, 
      pipeline_stageD_evaluate_jump_target_add_29_n190, 
      pipeline_stageD_evaluate_jump_target_add_29_n189, 
      pipeline_stageD_evaluate_jump_target_add_29_n188, 
      pipeline_stageD_evaluate_jump_target_add_29_n185, 
      pipeline_stageD_evaluate_jump_target_add_29_n184, 
      pipeline_stageD_evaluate_jump_target_add_29_n183, 
      pipeline_stageD_evaluate_jump_target_add_29_n182, 
      pipeline_stageD_evaluate_jump_target_add_29_n181, 
      pipeline_stageD_evaluate_jump_target_add_29_n180, 
      pipeline_stageD_evaluate_jump_target_add_29_n178, 
      pipeline_stageD_evaluate_jump_target_add_29_n177, 
      pipeline_stageD_evaluate_jump_target_add_29_n175, 
      pipeline_stageD_evaluate_jump_target_add_29_n174, 
      pipeline_stageD_evaluate_jump_target_add_29_n172, 
      pipeline_stageD_evaluate_jump_target_add_29_n171, 
      pipeline_stageD_evaluate_jump_target_add_29_n170, 
      pipeline_stageD_evaluate_jump_target_add_29_n169, 
      pipeline_stageD_evaluate_jump_target_add_29_n168, 
      pipeline_stageD_evaluate_jump_target_add_29_n165, 
      pipeline_stageD_evaluate_jump_target_add_29_n163, 
      pipeline_stageD_evaluate_jump_target_add_29_n160, 
      pipeline_stageD_evaluate_jump_target_add_29_n159, 
      pipeline_stageD_evaluate_jump_target_add_29_n157, 
      pipeline_stageD_evaluate_jump_target_add_29_n150, 
      pipeline_stageD_evaluate_jump_target_add_29_n149, 
      pipeline_stageD_evaluate_jump_target_add_29_n145, 
      pipeline_stageD_evaluate_jump_target_add_29_n144, 
      pipeline_stageD_evaluate_jump_target_add_29_n141, 
      pipeline_stageD_evaluate_jump_target_add_29_n139, 
      pipeline_stageD_evaluate_jump_target_add_29_n138, 
      pipeline_stageD_evaluate_jump_target_add_29_n135, 
      pipeline_stageD_evaluate_jump_target_add_29_n134, 
      pipeline_stageD_evaluate_jump_target_add_29_n133, 
      pipeline_stageD_evaluate_jump_target_add_29_n132, 
      pipeline_stageD_evaluate_jump_target_add_29_n129, 
      pipeline_stageD_evaluate_jump_target_add_29_n128, 
      pipeline_stageD_evaluate_jump_target_add_29_n126, n17018, n17019, n17020,
      n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028, n17029, 
      n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037, n17038, 
      n17039, n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047, 
      n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056, 
      n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065, 
      n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074, 
      n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083, 
      n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092, 
      n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101, 
      n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109, n17110, 
      n17111, n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119, 
      n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128, 
      n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137, 
      n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146, 
      n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155, 
      n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163, n17164, 
      n17165, n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173, 
      n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181, n17182, 
      n17183, n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191, 
      n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200, 
      n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209, 
      n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218, 
      n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227, 
      n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235, n17236, 
      n17237, n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245, 
      n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253, n17254, 
      n17255, n17256, n17257, n17258, n17259, n17260, n17261, n17262, n17263, 
      n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272, 
      n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281, 
      n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290, 
      n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299, 
      n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307, n17308, 
      n17309, n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317, 
      n17318, n17319, n17320, n17321, n17322, n17323, n17324, n17325, n17326, 
      n17327, n17328, n17329, n17330, n17331, n17332, n17333, n17334, n17335, 
      n17336, n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344, 
      n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353, 
      n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362, 
      n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371, 
      n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379, n17380, 
      n17381, n17382, n17383, n17384, n17385, n17386, n17387, n17388, n17389, 
      n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397, n17398, 
      n17399, n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407, 
      n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416, 
      n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425, 
      n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434, 
      n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443, 
      n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451, n17452, 
      n17453, n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461, 
      n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469, n17470, 
      n17471, n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479, 
      n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488, 
      n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497, 
      n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506, 
      n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515, 
      n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523, n17524, 
      n17525, n17526, n17527, n17528, n17529, n17530, n17531, n17532, n17533, 
      n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541, n17542, 
      n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17551, 
      n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560, 
      n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569, 
      n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578, 
      n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587, 
      n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595, n17596, 
      n17597, n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605, 
      n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614, 
      n17615, n17616, n17617, n17618, n17619, n17620, n17621, n17622, n17623, 
      n17624, n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632, 
      n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641, 
      n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650, 
      n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659, 
      n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667, n17668, 
      n17669, n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677, 
      n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686, 
      n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17695, 
      n17696, n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704, 
      n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713, 
      n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722, 
      n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731, 
      n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739, n17740, 
      n17741, n17742, n17743, n17744, net214675, net214676, net214677, 
      net214678, net214679, net214680, net214681, net214682, net214683, 
      net214684, net214685, net214686, net214687, net214688, net214689, 
      net214690, net214691, net214692, net214693, net214694, net214695, 
      net214696, net214697, net214698, net214699, net214700, net214701, 
      net214702, net214703, net214704, net214705, net214706, net214707, 
      net214708, net214709, net214710, net214711, net214712, net214713, 
      net214714, net214715, net214716, net214717, net214718, net214719, 
      net214720, net214721, net214722, net214723, net214724, net214725, 
      net214726, net214727, net214728, net214729, net214730, net214731, 
      net214732, net214733, net214734, net214735, net214736, net214737, 
      net214738, net214739, net214740, net214741, net214742, net214743, 
      net214744, net214745, net214746, net214747, net214748, net214749, 
      net214750, net214751, net214752, net214753, net214754, net214755, 
      net214756, net214757, net214758, net214759, net214760, net214761, 
      net214762, net214763, net214764, net214765, net214766, net214767, 
      net214768, net214769, net214770, net214771, net214772, net214773, 
      net214774, net214775, net214776, net214777, net214778, net214779, 
      net214780, net214781, net214782, net214783, net214784, net214785, 
      net214786, net214787, net214788, net214789, net214790, net214791, 
      net214792, net214793, net214794, net214795, net214796, net214797, 
      net214798, net214799, net214800, net214801, net214802, net214803, 
      net214804, net214805, net214806, net214807, net214808, net214809, 
      net214810, net214811, net214812, net214813, net214814, net214815, 
      net214816, net214817, net214818, net214819, net214820, net214821, 
      net214822, net214823, net214824, net214825 : std_logic;

begin
   
   DataMem_Mem_reg_7_31_inst : DLH_X1 port map( G => n13079, D => DataMem_N2159
                           , Q => DataMem_Mem_7_31_port);
   DataMem_Dataout_reg_31_inst : DLL_X1 port map( D => DataMem_N2254, GN => 
                           n17098, Q => DataMem_N2256);
   pipeline_MEMWB_Stage_Data_to_RF_reg_31_inst : DFF_X1 port map( D => 
                           pipeline_MEMWB_Stage_N42, CK => Clk, Q => 
                           pipeline_data_to_RF_from_WB_31_port, QN => n17425);
   pipeline_RegFile_DEC_WB_RegBank_reg_1_31_inst : DLH_X1 port map( G => n13172
                           , D => n13268, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_1_31_port);
   pipeline_IDEX_Stage_Reg1_out_IDEX_reg_31_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N133, CK => Clk, Q => n13966, QN
                           => net214825);
   pipeline_MEMWB_Stage_Data_to_RF_reg_0_inst : DFF_X1 port map( D => 
                           pipeline_MEMWB_Stage_N11, CK => Clk, Q => 
                           pipeline_data_to_RF_from_WB_0_port, QN => n17396);
   pipeline_RegFile_DEC_WB_RegBank_reg_1_0_inst : DLH_X1 port map( G => n17706,
                           D => n13175, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_1_0_port);
   pipeline_IDEX_Stage_Reg1_out_IDEX_reg_0_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N102, CK => Clk, Q => n13965, QN
                           => net214824);
   pipeline_MEMWB_Stage_Data_to_RF_reg_8_inst : DFF_X1 port map( D => 
                           pipeline_MEMWB_Stage_N19, CK => Clk, Q => 
                           pipeline_data_to_RF_from_WB_8_port, QN => n17394);
   pipeline_RegFile_DEC_WB_RegBank_reg_1_8_inst : DLH_X1 port map( G => n17706,
                           D => n13199, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_1_8_port);
   pipeline_IDEX_Stage_Reg1_out_IDEX_reg_8_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N110, CK => Clk, Q => n13964, QN
                           => net214823);
   pipeline_MEMWB_Stage_Data_to_RF_reg_24_inst : DFF_X1 port map( D => 
                           pipeline_MEMWB_Stage_N35, CK => Clk, Q => 
                           pipeline_data_to_RF_from_WB_24_port, QN => n17324);
   pipeline_RegFile_DEC_WB_RegBank_reg_1_24_inst : DLH_X1 port map( G => n13172
                           , D => n13247, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_1_24_port);
   pipeline_IDEX_Stage_Reg1_out_IDEX_reg_24_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N126, CK => Clk, Q => n13963, QN
                           => net214822);
   pipeline_MEMWB_Stage_Data_to_RF_reg_28_inst : DFF_X1 port map( D => 
                           pipeline_MEMWB_Stage_N39, CK => Clk, Q => 
                           pipeline_data_to_RF_from_WB_28_port, QN => n17312);
   pipeline_RegFile_DEC_WB_RegBank_reg_1_28_inst : DLH_X1 port map( G => n13172
                           , D => n13259, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_1_28_port);
   pipeline_IDEX_Stage_Reg1_out_IDEX_reg_28_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N130, CK => Clk, Q => n13962, QN
                           => net214821);
   pipeline_IFID_stage_Instr_out_IFID_reg_14_inst : DFF_X1 port map( D => n3992
                           , CK => Clk, Q => 
                           pipeline_stageD_offset_to_jump_temp_14_port, QN => 
                           n17445);
   pipeline_IDEX_Stage_Immediate_out_IDEX_reg_14_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N180, CK => Clk, Q => 
                           pipeline_immediate_to_exe_14_port, QN => net214820);
   pipeline_MEMWB_Stage_Data_to_RF_reg_14_inst : DFF_X1 port map( D => 
                           pipeline_MEMWB_Stage_N25, CK => Clk, Q => 
                           pipeline_data_to_RF_from_WB_14_port, QN => n17309);
   pipeline_RegFile_DEC_WB_RegBank_reg_1_14_inst : DLH_X1 port map( G => n13172
                           , D => n13217, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_1_14_port);
   pipeline_IDEX_Stage_Reg1_out_IDEX_reg_14_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N116, CK => Clk, Q => n13960, QN
                           => net214819);
   pipeline_MEMWB_Stage_Data_to_RF_reg_15_inst : DFF_X1 port map( D => 
                           pipeline_MEMWB_Stage_N26, CK => Clk, Q => 
                           pipeline_data_to_RF_from_WB_15_port, QN => n17364);
   pipeline_RegFile_DEC_WB_RegBank_reg_1_15_inst : DLH_X1 port map( G => n17706
                           , D => n13220, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_1_15_port);
   pipeline_IDEX_Stage_Reg1_out_IDEX_reg_15_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N117, CK => Clk, Q => n13959, QN
                           => net214818);
   pipeline_MEMWB_Stage_Data_to_RF_reg_13_inst : DFF_X1 port map( D => 
                           pipeline_MEMWB_Stage_N24, CK => Clk, Q => 
                           pipeline_data_to_RF_from_WB_13_port, QN => n17344);
   pipeline_RegFile_DEC_WB_RegBank_reg_1_13_inst : DLH_X1 port map( G => n13172
                           , D => n13214, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_1_13_port);
   pipeline_IDEX_Stage_Reg1_out_IDEX_reg_13_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N115, CK => Clk, Q => n13958, QN
                           => net214817);
   pipeline_MEMWB_Stage_Data_to_RF_reg_30_inst : DFF_X1 port map( D => 
                           pipeline_MEMWB_Stage_N41, CK => Clk, Q => 
                           pipeline_data_to_RF_from_WB_30_port, QN => n17362);
   pipeline_RegFile_DEC_WB_RegBank_reg_1_30_inst : DLH_X1 port map( G => n17706
                           , D => n13265, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_1_30_port);
   pipeline_IDEX_Stage_Reg1_out_IDEX_reg_30_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N132, CK => Clk, Q => n13957, QN
                           => net214816);
   pipeline_MEMWB_Stage_Data_to_RF_reg_29_inst : DFF_X1 port map( D => 
                           pipeline_MEMWB_Stage_N40, CK => Clk, Q => 
                           pipeline_data_to_RF_from_WB_29_port, QN => n17365);
   pipeline_RegFile_DEC_WB_RegBank_reg_1_29_inst : DLH_X1 port map( G => n17706
                           , D => n13262, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_1_29_port);
   pipeline_IDEX_Stage_Reg1_out_IDEX_reg_29_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N131, CK => Clk, Q => n13956, QN
                           => net214815);
   pipeline_MEMWB_Stage_Data_to_RF_reg_27_inst : DFF_X1 port map( D => 
                           pipeline_MEMWB_Stage_N38, CK => Clk, Q => 
                           pipeline_data_to_RF_from_WB_27_port, QN => n17325);
   pipeline_RegFile_DEC_WB_RegBank_reg_1_27_inst : DLH_X1 port map( G => n13172
                           , D => n13256, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_1_27_port);
   pipeline_IDEX_Stage_Reg1_out_IDEX_reg_27_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N129, CK => Clk, Q => n13955, QN
                           => net214814);
   pipeline_MEMWB_Stage_Data_to_RF_reg_26_inst : DFF_X1 port map( D => 
                           pipeline_MEMWB_Stage_N37, CK => Clk, Q => 
                           pipeline_data_to_RF_from_WB_26_port, QN => n17424);
   pipeline_RegFile_DEC_WB_RegBank_reg_1_26_inst : DLH_X1 port map( G => n13172
                           , D => n13253, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_1_26_port);
   pipeline_IDEX_Stage_Reg1_out_IDEX_reg_26_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N128, CK => Clk, Q => n13954, QN
                           => net214813);
   pipeline_MEMWB_Stage_Data_to_RF_reg_25_inst : DFF_X1 port map( D => 
                           pipeline_MEMWB_Stage_N36, CK => Clk, Q => 
                           pipeline_data_to_RF_from_WB_25_port, QN => n17427);
   pipeline_RegFile_DEC_WB_RegBank_reg_1_25_inst : DLH_X1 port map( G => n17706
                           , D => n13250, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_1_25_port);
   pipeline_IDEX_Stage_Reg1_out_IDEX_reg_25_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N127, CK => Clk, Q => n13953, QN
                           => net214812);
   pipeline_MEMWB_Stage_Data_to_RF_reg_23_inst : DFF_X1 port map( D => 
                           pipeline_MEMWB_Stage_N34, CK => Clk, Q => 
                           pipeline_data_to_RF_from_WB_23_port, QN => n17366);
   pipeline_RegFile_DEC_WB_RegBank_reg_1_23_inst : DLH_X1 port map( G => n17706
                           , D => n13244, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_1_23_port);
   pipeline_IDEX_Stage_Reg1_out_IDEX_reg_23_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N125, CK => Clk, Q => n13952, QN
                           => net214811);
   pipeline_MEMWB_Stage_Data_to_RF_reg_22_inst : DFF_X1 port map( D => 
                           pipeline_MEMWB_Stage_N33, CK => Clk, Q => 
                           pipeline_data_to_RF_from_WB_22_port, QN => n17311);
   pipeline_RegFile_DEC_WB_RegBank_reg_1_22_inst : DLH_X1 port map( G => n13172
                           , D => n13241, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_1_22_port);
   pipeline_IDEX_Stage_Reg1_out_IDEX_reg_22_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N124, CK => Clk, Q => n13951, QN
                           => net214810);
   pipeline_MEMWB_Stage_Data_to_RF_reg_21_inst : DFF_X1 port map( D => 
                           pipeline_MEMWB_Stage_N32, CK => Clk, Q => 
                           pipeline_data_to_RF_from_WB_21_port, QN => n17310);
   pipeline_RegFile_DEC_WB_RegBank_reg_1_21_inst : DLH_X1 port map( G => n13172
                           , D => n13238, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_1_21_port);
   pipeline_IDEX_Stage_Reg1_out_IDEX_reg_21_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N123, CK => Clk, Q => n13950, QN
                           => net214809);
   pipeline_MEMWB_Stage_Data_to_RF_reg_20_inst : DFF_X1 port map( D => 
                           pipeline_MEMWB_Stage_N31, CK => Clk, Q => 
                           pipeline_data_to_RF_from_WB_20_port, QN => n17322);
   pipeline_RegFile_DEC_WB_RegBank_reg_1_20_inst : DLH_X1 port map( G => n13172
                           , D => n13235, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_1_20_port);
   pipeline_IDEX_Stage_Reg1_out_IDEX_reg_20_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N122, CK => Clk, Q => n13949, QN
                           => net214808);
   pipeline_MEMWB_Stage_Data_to_RF_reg_19_inst : DFF_X1 port map( D => 
                           pipeline_MEMWB_Stage_N30, CK => Clk, Q => 
                           pipeline_data_to_RF_from_WB_19_port, QN => n17423);
   pipeline_RegFile_DEC_WB_RegBank_reg_1_19_inst : DLH_X1 port map( G => n17706
                           , D => n13232, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_1_19_port);
   pipeline_IDEX_Stage_Reg1_out_IDEX_reg_19_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N121, CK => Clk, Q => n13948, QN
                           => net214807);
   pipeline_MEMWB_Stage_Data_to_RF_reg_18_inst : DFF_X1 port map( D => 
                           pipeline_MEMWB_Stage_N29, CK => Clk, Q => 
                           pipeline_data_to_RF_from_WB_18_port, QN => n17363);
   pipeline_RegFile_DEC_WB_RegBank_reg_1_18_inst : DLH_X1 port map( G => n17706
                           , D => n13229, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_1_18_port);
   pipeline_IDEX_Stage_Reg1_out_IDEX_reg_18_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N120, CK => Clk, Q => n13947, QN
                           => net214806);
   pipeline_MEMWB_Stage_Data_to_RF_reg_17_inst : DFF_X1 port map( D => 
                           pipeline_MEMWB_Stage_N28, CK => Clk, Q => 
                           pipeline_data_to_RF_from_WB_17_port, QN => n17323);
   pipeline_RegFile_DEC_WB_RegBank_reg_1_17_inst : DLH_X1 port map( G => n13172
                           , D => n13226, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_1_17_port);
   pipeline_IDEX_Stage_Reg1_out_IDEX_reg_17_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N119, CK => Clk, Q => n13946, QN
                           => net214805);
   pipeline_MEMWB_Stage_Data_to_RF_reg_16_inst : DFF_X1 port map( D => 
                           pipeline_MEMWB_Stage_N27, CK => Clk, Q => 
                           pipeline_data_to_RF_from_WB_16_port, QN => n17426);
   pipeline_RegFile_DEC_WB_RegBank_reg_1_16_inst : DLH_X1 port map( G => n17706
                           , D => n13223, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_1_16_port);
   pipeline_stageF_PC_reg_PC_out_reg_16_inst : DFFR_X1 port map( D => n3991, CK
                           => Clk, RN => n17704, Q => n13945, QN => n7711);
   pipeline_IFID_stage_PC_out_IFID_reg_16_inst : DFF_X1 port map( D => n3990, 
                           CK => Clk, Q => pipeline_nextPC_IFID_DEC_16_port, QN
                           => n17461);
   pipeline_stageF_PC_reg_PC_out_reg_29_inst : DFFR_X1 port map( D => n3988, CK
                           => Clk, RN => n17704, Q => n13944, QN => n7709);
   pipeline_IFID_stage_Instr_out_IFID_reg_2_inst : DFF_X1 port map( D => n3985,
                           CK => Clk, Q => 
                           pipeline_stageD_offset_to_jump_temp_2_port, QN => 
                           n17404);
   pipeline_IFID_stage_Instr_out_IFID_reg_3_inst : DFF_X1 port map( D => n3984,
                           CK => Clk, Q => 
                           pipeline_stageD_offset_to_jump_temp_3_port, QN => 
                           n17410);
   pipeline_IFID_stage_Instr_out_IFID_reg_6_inst : DFF_X1 port map( D => n3981,
                           CK => Clk, Q => 
                           pipeline_stageD_offset_to_jump_temp_6_port, QN => 
                           n17361);
   pipeline_IFID_stage_Instr_out_IFID_reg_7_inst : DFF_X1 port map( D => n3980,
                           CK => Clk, Q => 
                           pipeline_stageD_offset_to_jump_temp_7_port, QN => 
                           n17437);
   pipeline_IFID_stage_Instr_out_IFID_reg_8_inst : DFF_X1 port map( D => n3979,
                           CK => Clk, Q => 
                           pipeline_stageD_offset_to_jump_temp_8_port, QN => 
                           n17428);
   pipeline_IFID_stage_Instr_out_IFID_reg_9_inst : DFF_X1 port map( D => n3978,
                           CK => Clk, Q => 
                           pipeline_stageD_offset_to_jump_temp_9_port, QN => 
                           n17432);
   pipeline_IFID_stage_Instr_out_IFID_reg_10_inst : DFF_X1 port map( D => n3977
                           , CK => Clk, Q => 
                           pipeline_stageD_offset_to_jump_temp_10_port, QN => 
                           n17440);
   pipeline_IFID_stage_Instr_out_IFID_reg_11_inst : DFF_X1 port map( D => n3976
                           , CK => Clk, Q => 
                           pipeline_stageD_offset_to_jump_temp_11_port, QN => 
                           n17433);
   pipeline_IFID_stage_Instr_out_IFID_reg_12_inst : DFF_X1 port map( D => n3975
                           , CK => Clk, Q => 
                           pipeline_stageD_offset_to_jump_temp_12_port, QN => 
                           n17444);
   pipeline_IFID_stage_Instr_out_IFID_reg_13_inst : DFF_X1 port map( D => n3974
                           , CK => Clk, Q => 
                           pipeline_stageD_offset_to_jump_temp_13_port, QN => 
                           n17434);
   pipeline_IFID_stage_Instr_out_IFID_reg_15_inst : DFF_X1 port map( D => n3973
                           , CK => Clk, Q => 
                           pipeline_stageD_offset_to_jump_temp_15_port, QN => 
                           n17431);
   pipeline_IFID_stage_Instr_out_IFID_reg_16_inst : DFF_X1 port map( D => n3972
                           , CK => Clk, Q => 
                           pipeline_stageD_offset_jump_sign_ext_16_port, QN => 
                           n17316);
   pipeline_IFID_stage_Instr_out_IFID_reg_17_inst : DFF_X1 port map( D => n3971
                           , CK => Clk, Q => 
                           pipeline_stageD_offset_jump_sign_ext_17_port, QN => 
                           n17329);
   pipeline_IFID_stage_Instr_out_IFID_reg_18_inst : DFF_X1 port map( D => n3970
                           , CK => Clk, Q => 
                           pipeline_stageD_offset_jump_sign_ext_18_port, QN => 
                           n17408);
   pipeline_IFID_stage_Instr_out_IFID_reg_19_inst : DFF_X1 port map( D => n3969
                           , CK => Clk, Q => 
                           pipeline_stageD_offset_jump_sign_ext_19_port, QN => 
                           n17349);
   pipeline_IFID_stage_Instr_out_IFID_reg_20_inst : DFF_X1 port map( D => n3968
                           , CK => Clk, Q => 
                           pipeline_stageD_offset_jump_sign_ext_20_port, QN => 
                           n17407);
   pipeline_IFID_stage_Instr_out_IFID_reg_26_inst : DFF_X1 port map( D => n3962
                           , CK => Clk, Q => pipeline_inst_IFID_DEC_26_port, QN
                           => n17409);
   pipeline_IFID_stage_Instr_out_IFID_reg_28_inst : DFF_X1 port map( D => n3960
                           , CK => Clk, Q => pipeline_inst_IFID_DEC_28_port, QN
                           => n17348);
   pipeline_IFID_stage_Instr_out_IFID_reg_30_inst : DFF_X1 port map( D => n3958
                           , CK => Clk, Q => pipeline_inst_IFID_DEC_30_port, QN
                           => n17347);
   pipeline_cu_pipeline_ALU_OPCODE_reg_2_inst : DLL_X1 port map( D => 
                           pipeline_cu_pipeline_N103, GN => Rst, Q => 
                           pipeline_EXE_controls_in_IDEX_3_port);
   pipeline_cu_pipeline_ALU_OPCODE_reg_3_inst : DLL_X1 port map( D => 
                           pipeline_cu_pipeline_N104, GN => Rst, Q => 
                           pipeline_EXE_controls_in_IDEX_4_port);
   pipeline_cu_pipeline_ALU_OPCODE_reg_5_inst : DLL_X1 port map( D => 
                           pipeline_cu_pipeline_N106, GN => Rst, Q => 
                           pipeline_EXE_controls_in_IDEX_6_port);
   pipeline_cu_pipeline_ALU_OPCODE_reg_0_inst : DLL_X1 port map( D => 
                           pipeline_cu_pipeline_N101, GN => Rst, Q => 
                           pipeline_EXE_controls_in_IDEX_1_port);
   pipeline_cu_pipeline_Reg_dst_reg : DLH_X1 port map( G => 
                           pipeline_cu_pipeline_N113, D => 
                           pipeline_cu_pipeline_N89, Q => 
                           pipeline_EXE_controls_in_IDEX_7_port);
   pipeline_cu_pipeline_Mem_to_reg_reg : DLH_X1 port map( G => 
                           pipeline_cu_pipeline_N107, D => 
                           pipeline_cu_pipeline_N108, Q => 
                           pipeline_WB_controls_in_IDEX_0_port);
   pipeline_cu_pipeline_ALU_OPCODE_reg_1_inst : DLL_X1 port map( D => 
                           pipeline_cu_pipeline_N102, GN => Rst, Q => 
                           pipeline_EXE_controls_in_IDEX_2_port);
   pipeline_cu_pipeline_Alu_src_reg : DLH_X1 port map( G => 
                           pipeline_cu_pipeline_N112, D => 
                           pipeline_cu_pipeline_N88, Q => 
                           pipeline_EXE_controls_in_IDEX_0_port);
   pipeline_cu_pipeline_isSigned_reg : DLH_X1 port map( G => 
                           pipeline_cu_pipeline_N109, D => 
                           pipeline_cu_pipeline_N110, Q => 
                           pipeline_EXE_controls_in_IDEX_8_port);
   pipeline_cu_pipeline_ALU_OPCODE_reg_4_inst : DLL_X1 port map( D => 
                           pipeline_cu_pipeline_N105, GN => Rst, Q => 
                           pipeline_EXE_controls_in_IDEX_5_port);
   pipeline_cu_hazard_stall_reg : DLH_X1 port map( G => pipeline_cu_hazard_N39,
                           D => pipeline_cu_hazard_N40, Q => pipeline_stall);
   pipeline_stageF_PC_reg_PC_out_tri_enable_reg_31_inst : DFFR_X1 port map( D 
                           => n3956, CK => Clk, RN => n17705, Q => 
                           pipeline_stageF_PC_reg_N0, QN => n17379);
   pipeline_stageF_PC_reg_PC_out_tri_enable_reg_29_inst : DFFR_X1 port map( D 
                           => n3955, CK => Clk, RN => n17704, Q => 
                           pipeline_stageF_PC_reg_N2, QN => n17494);
   pipeline_stageF_PC_reg_PC_out_tri_enable_reg_27_inst : DFFR_X1 port map( D 
                           => n3954, CK => Clk, RN => n17702, Q => 
                           pipeline_stageF_PC_reg_N4, QN => n17493);
   pipeline_stageF_PC_reg_PC_out_tri_enable_reg_25_inst : DFFR_X1 port map( D 
                           => n3953, CK => Clk, RN => n17705, Q => 
                           pipeline_stageF_PC_reg_N6, QN => n17492);
   pipeline_stageF_PC_reg_PC_out_tri_enable_reg_23_inst : DFFR_X1 port map( D 
                           => n3952, CK => Clk, RN => n17705, Q => 
                           pipeline_stageF_PC_reg_N8, QN => n17491);
   pipeline_stageF_PC_reg_PC_out_tri_enable_reg_21_inst : DFFR_X1 port map( D 
                           => n3951, CK => Clk, RN => n17703, Q => 
                           pipeline_stageF_PC_reg_N10, QN => n17490);
   pipeline_stageF_PC_reg_PC_out_tri_enable_reg_19_inst : DFFR_X1 port map( D 
                           => n3950, CK => Clk, RN => n17701, Q => 
                           pipeline_stageF_PC_reg_N12, QN => n17489);
   pipeline_stageF_PC_reg_PC_out_tri_enable_reg_17_inst : DFFR_X1 port map( D 
                           => n3949, CK => Clk, RN => n17705, Q => 
                           pipeline_stageF_PC_reg_N14, QN => n17488);
   pipeline_stageF_PC_reg_PC_out_tri_enable_reg_15_inst : DFFR_X1 port map( D 
                           => n3948, CK => Clk, RN => n17704, Q => 
                           pipeline_stageF_PC_reg_N16, QN => n17487);
   pipeline_stageF_PC_reg_PC_out_tri_enable_reg_13_inst : DFFR_X1 port map( D 
                           => n3947, CK => Clk, RN => n17704, Q => 
                           pipeline_stageF_PC_reg_N18, QN => n17486);
   pipeline_stageF_PC_reg_PC_out_tri_enable_reg_11_inst : DFFR_X1 port map( D 
                           => n3946, CK => Clk, RN => n17705, Q => 
                           pipeline_stageF_PC_reg_N20, QN => n17485);
   pipeline_stageF_PC_reg_PC_out_tri_enable_reg_9_inst : DFFR_X1 port map( D =>
                           n3945, CK => Clk, RN => n17705, Q => 
                           pipeline_stageF_PC_reg_N22, QN => n17378);
   pipeline_stageF_PC_reg_PC_out_tri_enable_reg_7_inst : DFFR_X1 port map( D =>
                           n3944, CK => Clk, RN => n17704, Q => 
                           pipeline_stageF_PC_reg_N24, QN => n17484);
   pipeline_stageF_PC_reg_PC_out_tri_enable_reg_5_inst : DFFR_X1 port map( D =>
                           n3943, CK => Clk, RN => n17705, Q => 
                           pipeline_stageF_PC_reg_N26, QN => n17483);
   pipeline_stageF_PC_reg_PC_out_tri_enable_reg_3_inst : DFFR_X1 port map( D =>
                           n3942, CK => Clk, RN => n17704, Q => 
                           pipeline_stageF_PC_reg_N28, QN => n17482);
   pipeline_stageF_PC_reg_PC_out_tri_enable_reg_1_inst : DFFR_X1 port map( D =>
                           n3941, CK => Clk, RN => n17705, Q => 
                           pipeline_stageF_PC_reg_N30, QN => n17377);
   pipeline_stageF_PC_reg_PC_out_tri_enable_reg_0_inst : DFFR_X1 port map( D =>
                           n3940, CK => Clk, RN => n17705, Q => 
                           pipeline_stageF_PC_reg_N31, QN => n17376);
   pipeline_stageF_PC_reg_PC_out_tri_enable_reg_2_inst : DFFR_X1 port map( D =>
                           n3939, CK => Clk, RN => n17704, Q => 
                           pipeline_stageF_PC_reg_N29, QN => n17481);
   pipeline_stageF_PC_reg_PC_out_tri_enable_reg_4_inst : DFFR_X1 port map( D =>
                           n3938, CK => Clk, RN => n17705, Q => 
                           pipeline_stageF_PC_reg_N27, QN => n17480);
   pipeline_stageF_PC_reg_PC_out_tri_enable_reg_6_inst : DFFR_X1 port map( D =>
                           n3937, CK => Clk, RN => n17704, Q => 
                           pipeline_stageF_PC_reg_N25, QN => n17479);
   pipeline_stageF_PC_reg_PC_out_tri_enable_reg_8_inst : DFFR_X1 port map( D =>
                           n3936, CK => Clk, RN => n17705, Q => 
                           pipeline_stageF_PC_reg_N23, QN => n17478);
   pipeline_stageF_PC_reg_PC_out_tri_enable_reg_10_inst : DFFR_X1 port map( D 
                           => n3935, CK => Clk, RN => n17705, Q => 
                           pipeline_stageF_PC_reg_N21, QN => n17375);
   pipeline_stageF_PC_reg_PC_out_tri_enable_reg_12_inst : DFFR_X1 port map( D 
                           => n3934, CK => Clk, RN => n17703, Q => 
                           pipeline_stageF_PC_reg_N19, QN => n17477);
   pipeline_stageF_PC_reg_PC_out_tri_enable_reg_14_inst : DFFR_X1 port map( D 
                           => n3933, CK => Clk, RN => n17702, Q => 
                           pipeline_stageF_PC_reg_N17, QN => n17476);
   pipeline_stageF_PC_reg_PC_out_tri_enable_reg_16_inst : DFFR_X1 port map( D 
                           => n3932, CK => Clk, RN => n17705, Q => 
                           pipeline_stageF_PC_reg_N15, QN => n17475);
   pipeline_stageF_PC_reg_PC_out_tri_enable_reg_18_inst : DFFR_X1 port map( D 
                           => n3931, CK => Clk, RN => n17704, Q => 
                           pipeline_stageF_PC_reg_N13, QN => n17474);
   pipeline_stageF_PC_reg_PC_out_tri_enable_reg_20_inst : DFFR_X1 port map( D 
                           => n3930, CK => Clk, RN => n17701, Q => 
                           pipeline_stageF_PC_reg_N11, QN => n17473);
   pipeline_stageF_PC_reg_PC_out_tri_enable_reg_22_inst : DFFR_X1 port map( D 
                           => n3929, CK => Clk, RN => n17705, Q => 
                           pipeline_stageF_PC_reg_N9, QN => n17374);
   pipeline_stageF_PC_reg_PC_out_tri_enable_reg_24_inst : DFFR_X1 port map( D 
                           => n3928, CK => Clk, RN => n17704, Q => 
                           pipeline_stageF_PC_reg_N7, QN => n17472);
   pipeline_stageF_PC_reg_PC_out_tri_enable_reg_26_inst : DFFR_X1 port map( D 
                           => n3927, CK => Clk, RN => n17705, Q => 
                           pipeline_stageF_PC_reg_N5, QN => n17373);
   pipeline_stageF_PC_reg_PC_out_tri_enable_reg_28_inst : DFFR_X1 port map( D 
                           => n3926, CK => Clk, RN => n17705, Q => 
                           pipeline_stageF_PC_reg_N3, QN => n17372);
   pipeline_stageF_PC_reg_PC_out_tri_enable_reg_30_inst : DFFR_X1 port map( D 
                           => n3925, CK => Clk, RN => n17705, Q => 
                           pipeline_stageF_PC_reg_N1, QN => n17371);
   pipeline_IDEX_Stage_MEM_controls_out_IDEX_reg_1_inst : DFF_X1 port map( D =>
                           pipeline_IDEX_Stage_N92, CK => Clk, Q => 
                           pipeline_MEM_controls_in_EXMEM_1_port, QN => 
                           net214804);
   pipeline_EXMEM_stage_MEM_controls_out_EXMEM_reg_1_inst : DFF_X1 port map( D 
                           => pipeline_EXMEM_stage_N6, CK => Clk, Q => 
                           pipeline_MEM_controls_in_MEM_1_port, QN => n17019);
   pipeline_IDEX_Stage_MEM_controls_out_IDEX_reg_0_inst : DFF_X1 port map( D =>
                           pipeline_IDEX_Stage_N91, CK => Clk, Q => n13942, QN 
                           => n17447);
   pipeline_EXMEM_stage_MEM_controls_out_EXMEM_reg_0_inst : DFF_X1 port map( D 
                           => pipeline_EXMEM_stage_N5, CK => Clk, Q => 
                           net214803, QN => n17020);
   pipeline_stageM_read_notWrite_reg : DLL_X1 port map( D => 
                           pipeline_MEM_controls_in_MEM_1_port, GN => n17155, Q
                           => read_notWrite);
   DataMem_Dataout_tri_enable_reg_31_inst : DLL_X1 port map( D => n17155, GN =>
                           n17098, Q => DataMem_N0);
   DataMem_Dataout_tri_enable_reg_29_inst : DLL_X1 port map( D => n12766, GN =>
                           n17098, Q => DataMem_N2);
   DataMem_Dataout_tri_enable_reg_27_inst : DLL_X1 port map( D => n12766, GN =>
                           n17098, Q => DataMem_N4);
   DataMem_Dataout_tri_enable_reg_25_inst : DLL_X1 port map( D => n17155, GN =>
                           n17098, Q => DataMem_N6);
   DataMem_Dataout_tri_enable_reg_23_inst : DLL_X1 port map( D => n17155, GN =>
                           n13055, Q => DataMem_N8);
   DataMem_Dataout_tri_enable_reg_21_inst : DLL_X1 port map( D => n12766, GN =>
                           n17098, Q => DataMem_N10);
   DataMem_Dataout_tri_enable_reg_19_inst : DLL_X1 port map( D => n17155, GN =>
                           n17098, Q => DataMem_N12);
   DataMem_Dataout_tri_enable_reg_17_inst : DLL_X1 port map( D => n12766, GN =>
                           n17098, Q => DataMem_N14);
   DataMem_Dataout_tri_enable_reg_15_inst : DLL_X1 port map( D => n12766, GN =>
                           n17098, Q => DataMem_N16);
   DataMem_Dataout_tri_enable_reg_13_inst : DLL_X1 port map( D => n17155, GN =>
                           n17098, Q => DataMem_N18);
   DataMem_Dataout_tri_enable_reg_11_inst : DLL_X1 port map( D => n12766, GN =>
                           n17098, Q => DataMem_N20);
   DataMem_Dataout_tri_enable_reg_9_inst : DLL_X1 port map( D => n17155, GN => 
                           n17098, Q => DataMem_N22);
   DataMem_Dataout_tri_enable_reg_7_inst : DLL_X1 port map( D => n17155, GN => 
                           n17098, Q => DataMem_N24);
   DataMem_Dataout_tri_enable_reg_5_inst : DLL_X1 port map( D => n12766, GN => 
                           n17098, Q => DataMem_N26);
   DataMem_Dataout_tri_enable_reg_3_inst : DLL_X1 port map( D => n17155, GN => 
                           n17098, Q => DataMem_N28);
   DataMem_Dataout_tri_enable_reg_1_inst : DLL_X1 port map( D => n12766, GN => 
                           n17098, Q => DataMem_N30);
   DataMem_Dataout_tri_enable_reg_0_inst : DLL_X1 port map( D => n17155, GN => 
                           n17098, Q => DataMem_N31);
   DataMem_Dataout_tri_enable_reg_2_inst : DLL_X1 port map( D => n12766, GN => 
                           n17098, Q => DataMem_N29);
   DataMem_Dataout_tri_enable_reg_4_inst : DLL_X1 port map( D => n17155, GN => 
                           n17098, Q => DataMem_N27);
   DataMem_Dataout_tri_enable_reg_6_inst : DLL_X1 port map( D => n17155, GN => 
                           n17098, Q => DataMem_N25);
   DataMem_Dataout_tri_enable_reg_8_inst : DLL_X1 port map( D => n12766, GN => 
                           n17098, Q => DataMem_N23);
   DataMem_Dataout_tri_enable_reg_10_inst : DLL_X1 port map( D => n17155, GN =>
                           n17098, Q => DataMem_N21);
   DataMem_Dataout_tri_enable_reg_12_inst : DLL_X1 port map( D => n12766, GN =>
                           n17098, Q => DataMem_N19);
   DataMem_Dataout_tri_enable_reg_14_inst : DLL_X1 port map( D => n12766, GN =>
                           n17098, Q => DataMem_N17);
   DataMem_Dataout_tri_enable_reg_16_inst : DLL_X1 port map( D => n17155, GN =>
                           n17098, Q => DataMem_N15);
   DataMem_Dataout_tri_enable_reg_18_inst : DLL_X1 port map( D => n17155, GN =>
                           n17098, Q => DataMem_N13);
   DataMem_Dataout_tri_enable_reg_20_inst : DLL_X1 port map( D => n17155, GN =>
                           n17098, Q => DataMem_N11);
   DataMem_Dataout_tri_enable_reg_22_inst : DLL_X1 port map( D => n17155, GN =>
                           n17098, Q => DataMem_N9);
   DataMem_Dataout_tri_enable_reg_24_inst : DLL_X1 port map( D => n12766, GN =>
                           n17098, Q => DataMem_N7);
   DataMem_Dataout_tri_enable_reg_26_inst : DLL_X1 port map( D => n12766, GN =>
                           n17098, Q => DataMem_N5);
   DataMem_Dataout_tri_enable_reg_28_inst : DLL_X1 port map( D => n12766, GN =>
                           n17098, Q => DataMem_N3);
   DataMem_Dataout_tri_enable_reg_30_inst : DLL_X1 port map( D => n17155, GN =>
                           n17098, Q => DataMem_N1);
   pipeline_IDEX_Stage_WB_controls_out_IDEX_reg_1_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N90, CK => Clk, Q => 
                           pipeline_WB_controls_in_EXMEM_1_port, QN => n17449);
   pipeline_EXMEM_stage_WB_controls_out_EXMEM_reg_1_inst : DFF_X1 port map( D 
                           => pipeline_EXMEM_stage_N4, CK => Clk, Q => 
                           pipeline_WB_controls_in_MEMWB_1_port, QN => n17387);
   pipeline_MEMWB_Stage_writeback_reg : DFF_X1 port map( D => 
                           pipeline_MEMWB_Stage_N10, CK => Clk, Q => net214802,
                           QN => n13940);
   pipeline_IDEX_Stage_EXE_controls_out_IDEX_reg_8_inst : DFF_X1 port map( D =>
                           pipeline_IDEX_Stage_N101, CK => Clk, Q => n13939, QN
                           => net214801);
   pipeline_stageF_PC_reg_PC_out_reg_31_inst : DFFR_X1 port map( D => n3924, CK
                           => Clk, RN => n17705, Q => n13938, QN => n7676);
   pipeline_IFID_stage_PC_out_IFID_reg_31_inst : DFF_X1 port map( D => n3923, 
                           CK => Clk, Q => n13937, QN => n17527);
   pipeline_IDEX_Stage_EXE_controls_out_IDEX_reg_6_inst : DFF_X1 port map( D =>
                           pipeline_IDEX_Stage_N99, CK => Clk, Q => 
                           pipeline_EXE_controls_in_EXEcute_6_port, QN => 
                           n17421);
   pipeline_IDEX_Stage_EXE_controls_out_IDEX_reg_5_inst : DFF_X1 port map( D =>
                           pipeline_IDEX_Stage_N98, CK => Clk, Q => 
                           pipeline_EXE_controls_in_EXEcute_5_port, QN => 
                           net214800);
   pipeline_IDEX_Stage_EXE_controls_out_IDEX_reg_4_inst : DFF_X1 port map( D =>
                           pipeline_IDEX_Stage_N97, CK => Clk, Q => 
                           pipeline_EXE_controls_in_EXEcute_4_port, QN => 
                           net214799);
   pipeline_IDEX_Stage_EXE_controls_out_IDEX_reg_3_inst : DFF_X1 port map( D =>
                           pipeline_IDEX_Stage_N96, CK => Clk, Q => 
                           pipeline_EXE_controls_in_EXEcute_3_port, QN => 
                           n17411);
   pipeline_IDEX_Stage_EXE_controls_out_IDEX_reg_2_inst : DFF_X1 port map( D =>
                           pipeline_IDEX_Stage_N95, CK => Clk, Q => 
                           pipeline_EXE_controls_in_EXEcute_2_port, QN => 
                           n17405);
   pipeline_IDEX_Stage_WB_controls_out_IDEX_reg_0_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N89, CK => Clk, Q => n13936, QN 
                           => net214798);
   pipeline_EXMEM_stage_WB_controls_out_EXMEM_reg_0_inst : DFF_X1 port map( D 
                           => pipeline_EXMEM_stage_N3, CK => Clk, Q => 
                           pipeline_WB_controls_in_MEMWB_0_port, QN => 
                           net214797);
   pipeline_IDEX_Stage_RegDst_2_Addr_out_IDEX_reg_4_inst : DFF_X1 port map( D 
                           => pipeline_IDEX_Stage_N217, CK => Clk, Q => n13934,
                           QN => net214796);
   pipeline_IDEX_Stage_RegDst_2_Addr_out_IDEX_reg_3_inst : DFF_X1 port map( D 
                           => pipeline_IDEX_Stage_N216, CK => Clk, Q => n13933,
                           QN => net214795);
   pipeline_IDEX_Stage_RegDst_2_Addr_out_IDEX_reg_2_inst : DFF_X1 port map( D 
                           => pipeline_IDEX_Stage_N215, CK => Clk, Q => n13932,
                           QN => net214794);
   pipeline_IDEX_Stage_RegDst_2_Addr_out_IDEX_reg_1_inst : DFF_X1 port map( D 
                           => pipeline_IDEX_Stage_N214, CK => Clk, Q => n13931,
                           QN => net214793);
   pipeline_IDEX_Stage_RegDst_2_Addr_out_IDEX_reg_0_inst : DFF_X1 port map( D 
                           => pipeline_IDEX_Stage_N213, CK => Clk, Q => n13930,
                           QN => net214792);
   pipeline_IDEX_Stage_RegDst_1_Addr_out_IDEX_reg_4_inst : DFF_X1 port map( D 
                           => pipeline_IDEX_Stage_N212, CK => Clk, Q => n13929,
                           QN => net214791);
   pipeline_IDEX_Stage_RegDst_1_Addr_out_IDEX_reg_3_inst : DFF_X1 port map( D 
                           => pipeline_IDEX_Stage_N211, CK => Clk, Q => n13928,
                           QN => net214790);
   pipeline_IDEX_Stage_RegDst_1_Addr_out_IDEX_reg_2_inst : DFF_X1 port map( D 
                           => pipeline_IDEX_Stage_N210, CK => Clk, Q => n13927,
                           QN => net214789);
   pipeline_IDEX_Stage_RegDst_1_Addr_out_IDEX_reg_1_inst : DFF_X1 port map( D 
                           => pipeline_IDEX_Stage_N209, CK => Clk, Q => n13926,
                           QN => net214788);
   pipeline_IDEX_Stage_RegDst_1_Addr_out_IDEX_reg_0_inst : DFF_X1 port map( D 
                           => pipeline_IDEX_Stage_N208, CK => Clk, Q => n13925,
                           QN => net214787);
   pipeline_IDEX_Stage_Immediate_out_IDEX_reg_2_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N168, CK => Clk, Q => 
                           pipeline_immediate_to_exe_2_port, QN => net214786);
   pipeline_IDEX_Stage_Reg2_Addr_out_IDEX_reg_3_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N206, CK => Clk, Q => 
                           pipeline_Reg2_Addr_to_exe_3_port, QN => net214785);
   pipeline_IDEX_Stage_Reg2_Addr_out_IDEX_reg_2_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N205, CK => Clk, Q => 
                           pipeline_Reg2_Addr_to_exe_2_port, QN => n17403);
   pipeline_IDEX_Stage_Reg2_Addr_out_IDEX_reg_0_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N203, CK => Clk, Q => 
                           pipeline_Reg2_Addr_to_exe_0_port, QN => net214784);
   pipeline_IDEX_Stage_Reg1_Addr_out_IDEX_reg_4_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N202, CK => Clk, Q => 
                           pipeline_Reg1_Addr_to_exe_4_port, QN => n17399);
   pipeline_IDEX_Stage_Reg1_Addr_out_IDEX_reg_3_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N201, CK => Clk, Q => 
                           pipeline_Reg1_Addr_to_exe_3_port, QN => net214783);
   pipeline_IDEX_Stage_Reg1_Addr_out_IDEX_reg_2_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N200, CK => Clk, Q => 
                           pipeline_Reg1_Addr_to_exe_2_port, QN => n17401);
   pipeline_IDEX_Stage_Reg1_Addr_out_IDEX_reg_1_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N199, CK => Clk, Q => 
                           pipeline_Reg1_Addr_to_exe_1_port, QN => net214782);
   pipeline_IDEX_Stage_Immediate_out_IDEX_reg_15_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N181, CK => Clk, Q => 
                           pipeline_immediate_to_exe_15_port, QN => net214781);
   pipeline_IDEX_Stage_Immediate_out_IDEX_reg_13_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N179, CK => Clk, Q => 
                           pipeline_immediate_to_exe_13_port, QN => net214780);
   pipeline_IDEX_Stage_Immediate_out_IDEX_reg_12_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N178, CK => Clk, Q => 
                           pipeline_immediate_to_exe_12_port, QN => net214779);
   pipeline_IDEX_Stage_Immediate_out_IDEX_reg_11_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N177, CK => Clk, Q => 
                           pipeline_immediate_to_exe_11_port, QN => net214778);
   pipeline_IDEX_Stage_Immediate_out_IDEX_reg_9_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N175, CK => Clk, Q => 
                           pipeline_immediate_to_exe_9_port, QN => net214777);
   pipeline_IDEX_Stage_Immediate_out_IDEX_reg_8_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N174, CK => Clk, Q => 
                           pipeline_immediate_to_exe_8_port, QN => net214776);
   pipeline_IDEX_Stage_Immediate_out_IDEX_reg_7_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N173, CK => Clk, Q => 
                           pipeline_immediate_to_exe_7_port, QN => net214775);
   pipeline_IDEX_Stage_Immediate_out_IDEX_reg_31_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N197, CK => Clk, Q => 
                           pipeline_immediate_to_exe_31_port, QN => net214774);
   pipeline_IDEX_Stage_Immediate_out_IDEX_reg_29_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N197, CK => Clk, Q => 
                           pipeline_immediate_to_exe_29_port, QN => net214773);
   pipeline_IDEX_Stage_Immediate_out_IDEX_reg_27_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N197, CK => Clk, Q => 
                           pipeline_immediate_to_exe_27_port, QN => net214772);
   pipeline_IDEX_Stage_Immediate_out_IDEX_reg_25_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N197, CK => Clk, Q => 
                           pipeline_immediate_to_exe_25_port, QN => net214771);
   pipeline_IDEX_Stage_Immediate_out_IDEX_reg_23_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N197, CK => Clk, Q => 
                           pipeline_immediate_to_exe_23_port, QN => net214770);
   pipeline_IDEX_Stage_Immediate_out_IDEX_reg_21_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N197, CK => Clk, Q => 
                           pipeline_immediate_to_exe_21_port, QN => net214769);
   pipeline_IDEX_Stage_Immediate_out_IDEX_reg_19_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N197, CK => Clk, Q => 
                           pipeline_immediate_to_exe_19_port, QN => net214768);
   pipeline_IDEX_Stage_Immediate_out_IDEX_reg_17_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N197, CK => Clk, Q => 
                           pipeline_immediate_to_exe_17_port, QN => net214767);
   pipeline_IDEX_Stage_Immediate_out_IDEX_reg_16_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N197, CK => Clk, Q => 
                           pipeline_immediate_to_exe_16_port, QN => net214766);
   pipeline_IDEX_Stage_Immediate_out_IDEX_reg_18_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N197, CK => Clk, Q => 
                           pipeline_immediate_to_exe_18_port, QN => net214765);
   pipeline_IDEX_Stage_Immediate_out_IDEX_reg_20_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N197, CK => Clk, Q => 
                           pipeline_immediate_to_exe_20_port, QN => net214764);
   pipeline_IDEX_Stage_Immediate_out_IDEX_reg_22_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N197, CK => Clk, Q => 
                           pipeline_immediate_to_exe_22_port, QN => net214763);
   pipeline_IDEX_Stage_Immediate_out_IDEX_reg_24_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N197, CK => Clk, Q => 
                           pipeline_immediate_to_exe_24_port, QN => net214762);
   pipeline_IDEX_Stage_Immediate_out_IDEX_reg_26_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N197, CK => Clk, Q => 
                           pipeline_immediate_to_exe_26_port, QN => net214761);
   pipeline_IDEX_Stage_Immediate_out_IDEX_reg_28_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N197, CK => Clk, Q => 
                           pipeline_immediate_to_exe_28_port, QN => net214760);
   pipeline_IDEX_Stage_Immediate_out_IDEX_reg_30_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N197, CK => Clk, Q => 
                           pipeline_immediate_to_exe_30_port, QN => net214759);
   pipeline_IDEX_Stage_Immediate_out_IDEX_reg_10_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N176, CK => Clk, Q => 
                           pipeline_immediate_to_exe_10_port, QN => net214758);
   pipeline_IDEX_Stage_Immediate_out_IDEX_reg_6_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N172, CK => Clk, Q => 
                           pipeline_immediate_to_exe_6_port, QN => net214757);
   pipeline_IDEX_Stage_Immediate_out_IDEX_reg_5_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N171, CK => Clk, Q => 
                           pipeline_immediate_to_exe_5_port, QN => net214756);
   pipeline_IDEX_Stage_Immediate_out_IDEX_reg_4_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N170, CK => Clk, Q => 
                           pipeline_immediate_to_exe_4_port, QN => net214755);
   pipeline_IDEX_Stage_Immediate_out_IDEX_reg_3_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N169, CK => Clk, Q => 
                           pipeline_immediate_to_exe_3_port, QN => net214754);
   pipeline_IDEX_Stage_Immediate_out_IDEX_reg_1_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N167, CK => Clk, Q => 
                           pipeline_immediate_to_exe_1_port, QN => net214753);
   pipeline_IDEX_Stage_Immediate_out_IDEX_reg_0_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N166, CK => Clk, Q => net214752,
                           QN => n17400);
   pipeline_IDEX_Stage_EXE_controls_out_IDEX_reg_7_inst : DFF_X1 port map( D =>
                           pipeline_IDEX_Stage_N100, CK => Clk, Q => 
                           pipeline_EXE_controls_in_EXEcute_7_port, QN => 
                           n17430);
   pipeline_MEMWB_Stage_RegDst_Addr_out_MEMWB_reg_3_inst : DFF_X1 port map( D 
                           => pipeline_MEMWB_Stage_N46, CK => Clk, Q => 
                           pipeline_RegDst_to_WB_3_port, QN => n17385);
   pipeline_RegFile_DEC_WB_RegBank_reg_2_31_inst : DLH_X1 port map( G => n13169
                           , D => n13268, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_2_31_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_2_29_inst : DLH_X1 port map( G => n17707
                           , D => n13262, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_2_29_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_2_27_inst : DLH_X1 port map( G => n13169
                           , D => n13256, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_2_27_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_2_25_inst : DLH_X1 port map( G => n17707
                           , D => n13250, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_2_25_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_2_23_inst : DLH_X1 port map( G => n17707
                           , D => n13244, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_2_23_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_2_21_inst : DLH_X1 port map( G => n13169
                           , D => n13238, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_2_21_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_2_19_inst : DLH_X1 port map( G => n17707
                           , D => n13232, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_2_19_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_2_17_inst : DLH_X1 port map( G => n13169
                           , D => n13226, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_2_17_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_2_15_inst : DLH_X1 port map( G => n17707
                           , D => n13220, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_2_15_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_2_13_inst : DLH_X1 port map( G => n13169
                           , D => n13214, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_2_13_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_2_0_inst : DLH_X1 port map( G => n17707,
                           D => n13175, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_2_0_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_2_8_inst : DLH_X1 port map( G => n17707,
                           D => n13199, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_2_8_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_2_14_inst : DLH_X1 port map( G => n13169
                           , D => n13217, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_2_14_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_2_16_inst : DLH_X1 port map( G => n17707
                           , D => n13223, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_2_16_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_2_18_inst : DLH_X1 port map( G => n17707
                           , D => n13229, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_2_18_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_2_20_inst : DLH_X1 port map( G => n13169
                           , D => n13235, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_2_20_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_2_22_inst : DLH_X1 port map( G => n13169
                           , D => n13241, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_2_22_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_2_24_inst : DLH_X1 port map( G => n13169
                           , D => n13247, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_2_24_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_2_26_inst : DLH_X1 port map( G => n13169
                           , D => n13253, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_2_26_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_2_28_inst : DLH_X1 port map( G => n13169
                           , D => n13259, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_2_28_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_2_30_inst : DLH_X1 port map( G => n17707
                           , D => n13265, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_2_30_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_3_31_inst : DLH_X1 port map( G => n17708
                           , D => n13268, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_3_31_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_3_29_inst : DLH_X1 port map( G => n17708
                           , D => n13262, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_3_29_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_3_27_inst : DLH_X1 port map( G => n13166
                           , D => n13256, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_3_27_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_3_25_inst : DLH_X1 port map( G => n17708
                           , D => n13250, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_3_25_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_3_23_inst : DLH_X1 port map( G => n13166
                           , D => n13244, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_3_23_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_3_21_inst : DLH_X1 port map( G => n13166
                           , D => n13238, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_3_21_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_3_19_inst : DLH_X1 port map( G => n17708
                           , D => n13232, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_3_19_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_3_17_inst : DLH_X1 port map( G => n13166
                           , D => n13226, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_3_17_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_3_15_inst : DLH_X1 port map( G => n17708
                           , D => n13220, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_3_15_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_3_13_inst : DLH_X1 port map( G => n13166
                           , D => n13214, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_3_13_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_3_0_inst : DLH_X1 port map( G => n17708,
                           D => n13175, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_3_0_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_3_8_inst : DLH_X1 port map( G => n17708,
                           D => n13199, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_3_8_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_3_14_inst : DLH_X1 port map( G => n13166
                           , D => n13217, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_3_14_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_3_16_inst : DLH_X1 port map( G => n17708
                           , D => n13223, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_3_16_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_3_18_inst : DLH_X1 port map( G => n17708
                           , D => n13229, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_3_18_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_3_20_inst : DLH_X1 port map( G => n13166
                           , D => n13235, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_3_20_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_3_22_inst : DLH_X1 port map( G => n13166
                           , D => n13241, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_3_22_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_3_24_inst : DLH_X1 port map( G => n13166
                           , D => n13247, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_3_24_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_3_26_inst : DLH_X1 port map( G => n13166
                           , D => n13253, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_3_26_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_3_28_inst : DLH_X1 port map( G => n13166
                           , D => n13259, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_3_28_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_3_30_inst : DLH_X1 port map( G => n17708
                           , D => n13265, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_3_30_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_4_31_inst : DLH_X1 port map( G => n13163
                           , D => n13268, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_4_31_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_4_29_inst : DLH_X1 port map( G => n17709
                           , D => n13262, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_4_29_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_4_27_inst : DLH_X1 port map( G => n13163
                           , D => n13256, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_4_27_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_4_25_inst : DLH_X1 port map( G => n17709
                           , D => n13250, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_4_25_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_4_23_inst : DLH_X1 port map( G => n17709
                           , D => n13244, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_4_23_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_4_21_inst : DLH_X1 port map( G => n13163
                           , D => n13238, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_4_21_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_4_19_inst : DLH_X1 port map( G => n17709
                           , D => n13232, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_4_19_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_4_17_inst : DLH_X1 port map( G => n13163
                           , D => n13226, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_4_17_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_4_15_inst : DLH_X1 port map( G => n17709
                           , D => n13220, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_4_15_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_4_13_inst : DLH_X1 port map( G => n13163
                           , D => n13214, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_4_13_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_4_0_inst : DLH_X1 port map( G => n17709,
                           D => n13175, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_4_0_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_4_8_inst : DLH_X1 port map( G => n17709,
                           D => n13199, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_4_8_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_4_14_inst : DLH_X1 port map( G => n13163
                           , D => n13217, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_4_14_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_4_16_inst : DLH_X1 port map( G => n17709
                           , D => n13223, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_4_16_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_4_18_inst : DLH_X1 port map( G => n17709
                           , D => n13229, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_4_18_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_4_20_inst : DLH_X1 port map( G => n13163
                           , D => n13235, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_4_20_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_4_22_inst : DLH_X1 port map( G => n13163
                           , D => n13241, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_4_22_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_4_24_inst : DLH_X1 port map( G => n13163
                           , D => n13247, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_4_24_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_4_26_inst : DLH_X1 port map( G => n13163
                           , D => n13253, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_4_26_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_4_28_inst : DLH_X1 port map( G => n13163
                           , D => n13259, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_4_28_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_4_30_inst : DLH_X1 port map( G => n17709
                           , D => n13265, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_4_30_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_5_31_inst : DLH_X1 port map( G => n13160
                           , D => n13268, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_5_31_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_5_29_inst : DLH_X1 port map( G => n17710
                           , D => n13262, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_5_29_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_5_27_inst : DLH_X1 port map( G => n13160
                           , D => n13256, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_5_27_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_5_25_inst : DLH_X1 port map( G => n17710
                           , D => n13250, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_5_25_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_5_23_inst : DLH_X1 port map( G => n17710
                           , D => n13244, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_5_23_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_5_21_inst : DLH_X1 port map( G => n13160
                           , D => n13238, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_5_21_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_5_19_inst : DLH_X1 port map( G => n17710
                           , D => n13232, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_5_19_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_5_17_inst : DLH_X1 port map( G => n13160
                           , D => n13226, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_5_17_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_5_15_inst : DLH_X1 port map( G => n17710
                           , D => n13220, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_5_15_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_5_13_inst : DLH_X1 port map( G => n13160
                           , D => n13214, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_5_13_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_5_0_inst : DLH_X1 port map( G => n17710,
                           D => n13175, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_5_0_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_5_8_inst : DLH_X1 port map( G => n17710,
                           D => n13199, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_5_8_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_5_14_inst : DLH_X1 port map( G => n13160
                           , D => n13217, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_5_14_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_5_16_inst : DLH_X1 port map( G => n17710
                           , D => n13223, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_5_16_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_5_18_inst : DLH_X1 port map( G => n17710
                           , D => n13229, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_5_18_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_5_20_inst : DLH_X1 port map( G => n13160
                           , D => n13235, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_5_20_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_5_22_inst : DLH_X1 port map( G => n13160
                           , D => n13241, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_5_22_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_5_24_inst : DLH_X1 port map( G => n13160
                           , D => n13247, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_5_24_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_5_26_inst : DLH_X1 port map( G => n13160
                           , D => n13253, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_5_26_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_5_28_inst : DLH_X1 port map( G => n13160
                           , D => n13259, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_5_28_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_5_30_inst : DLH_X1 port map( G => n17710
                           , D => n13265, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_5_30_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_6_31_inst : DLH_X1 port map( G => n13157
                           , D => n13268, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_6_31_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_6_29_inst : DLH_X1 port map( G => n17711
                           , D => n13262, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_6_29_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_6_27_inst : DLH_X1 port map( G => n13157
                           , D => n13256, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_6_27_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_6_25_inst : DLH_X1 port map( G => n17711
                           , D => n13250, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_6_25_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_6_23_inst : DLH_X1 port map( G => n17711
                           , D => n13244, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_6_23_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_6_21_inst : DLH_X1 port map( G => n13157
                           , D => n13238, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_6_21_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_6_19_inst : DLH_X1 port map( G => n17711
                           , D => n13232, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_6_19_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_6_17_inst : DLH_X1 port map( G => n13157
                           , D => n13226, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_6_17_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_6_15_inst : DLH_X1 port map( G => n17711
                           , D => n13220, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_6_15_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_6_13_inst : DLH_X1 port map( G => n13157
                           , D => n13214, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_6_13_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_6_0_inst : DLH_X1 port map( G => n17711,
                           D => n13175, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_6_0_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_6_8_inst : DLH_X1 port map( G => n17711,
                           D => n13199, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_6_8_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_6_14_inst : DLH_X1 port map( G => n13157
                           , D => n13217, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_6_14_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_6_16_inst : DLH_X1 port map( G => n17711
                           , D => n13223, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_6_16_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_6_18_inst : DLH_X1 port map( G => n17711
                           , D => n13229, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_6_18_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_6_20_inst : DLH_X1 port map( G => n13157
                           , D => n13235, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_6_20_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_6_22_inst : DLH_X1 port map( G => n13157
                           , D => n13241, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_6_22_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_6_24_inst : DLH_X1 port map( G => n13157
                           , D => n13247, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_6_24_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_6_26_inst : DLH_X1 port map( G => n13157
                           , D => n13253, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_6_26_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_6_28_inst : DLH_X1 port map( G => n13157
                           , D => n13259, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_6_28_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_6_30_inst : DLH_X1 port map( G => n17711
                           , D => n13265, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_6_30_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_7_31_inst : DLH_X1 port map( G => n13154
                           , D => n13268, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_7_31_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_7_29_inst : DLH_X1 port map( G => n17712
                           , D => n13262, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_7_29_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_7_27_inst : DLH_X1 port map( G => n13154
                           , D => n13256, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_7_27_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_7_25_inst : DLH_X1 port map( G => n17712
                           , D => n13250, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_7_25_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_7_23_inst : DLH_X1 port map( G => n17712
                           , D => n13244, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_7_23_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_7_21_inst : DLH_X1 port map( G => n13154
                           , D => n13238, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_7_21_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_7_19_inst : DLH_X1 port map( G => n17712
                           , D => n13232, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_7_19_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_7_17_inst : DLH_X1 port map( G => n13154
                           , D => n13226, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_7_17_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_7_15_inst : DLH_X1 port map( G => n17712
                           , D => n13220, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_7_15_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_7_13_inst : DLH_X1 port map( G => n13154
                           , D => n13214, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_7_13_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_7_0_inst : DLH_X1 port map( G => n17712,
                           D => n13175, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_7_0_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_7_8_inst : DLH_X1 port map( G => n17712,
                           D => n13199, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_7_8_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_7_14_inst : DLH_X1 port map( G => n13154
                           , D => n13217, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_7_14_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_7_16_inst : DLH_X1 port map( G => n17712
                           , D => n13223, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_7_16_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_7_18_inst : DLH_X1 port map( G => n17712
                           , D => n13229, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_7_18_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_7_20_inst : DLH_X1 port map( G => n13154
                           , D => n13235, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_7_20_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_7_22_inst : DLH_X1 port map( G => n13154
                           , D => n13241, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_7_22_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_7_24_inst : DLH_X1 port map( G => n13154
                           , D => n13247, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_7_24_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_7_26_inst : DLH_X1 port map( G => n13154
                           , D => n13253, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_7_26_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_7_28_inst : DLH_X1 port map( G => n13154
                           , D => n13259, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_7_28_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_7_30_inst : DLH_X1 port map( G => n17712
                           , D => n13265, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_7_30_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_8_31_inst : DLH_X1 port map( G => n13151
                           , D => n13268, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_8_31_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_8_29_inst : DLH_X1 port map( G => n17713
                           , D => n13262, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_8_29_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_8_27_inst : DLH_X1 port map( G => n13151
                           , D => n13256, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_8_27_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_8_25_inst : DLH_X1 port map( G => n17713
                           , D => n13250, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_8_25_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_8_23_inst : DLH_X1 port map( G => n17713
                           , D => n13244, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_8_23_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_8_21_inst : DLH_X1 port map( G => n13151
                           , D => n13238, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_8_21_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_8_19_inst : DLH_X1 port map( G => n17713
                           , D => n13232, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_8_19_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_8_17_inst : DLH_X1 port map( G => n13151
                           , D => n13226, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_8_17_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_8_15_inst : DLH_X1 port map( G => n17713
                           , D => n13220, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_8_15_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_8_13_inst : DLH_X1 port map( G => n13151
                           , D => n13214, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_8_13_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_8_0_inst : DLH_X1 port map( G => n17713,
                           D => n13175, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_8_0_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_8_8_inst : DLH_X1 port map( G => n17713,
                           D => n13199, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_8_8_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_8_14_inst : DLH_X1 port map( G => n13151
                           , D => n13217, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_8_14_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_8_16_inst : DLH_X1 port map( G => n17713
                           , D => n13223, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_8_16_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_8_18_inst : DLH_X1 port map( G => n17713
                           , D => n13229, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_8_18_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_8_20_inst : DLH_X1 port map( G => n13151
                           , D => n13235, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_8_20_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_8_22_inst : DLH_X1 port map( G => n13151
                           , D => n13241, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_8_22_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_8_24_inst : DLH_X1 port map( G => n13151
                           , D => n13247, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_8_24_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_8_26_inst : DLH_X1 port map( G => n13151
                           , D => n13253, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_8_26_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_8_28_inst : DLH_X1 port map( G => n13151
                           , D => n13259, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_8_28_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_8_30_inst : DLH_X1 port map( G => n17713
                           , D => n13265, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_8_30_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_9_31_inst : DLH_X1 port map( G => n13148
                           , D => n13268, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_9_31_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_9_29_inst : DLH_X1 port map( G => n17714
                           , D => n13262, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_9_29_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_9_27_inst : DLH_X1 port map( G => n13148
                           , D => n13256, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_9_27_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_9_25_inst : DLH_X1 port map( G => n17714
                           , D => n13250, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_9_25_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_9_23_inst : DLH_X1 port map( G => n17714
                           , D => n13244, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_9_23_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_9_21_inst : DLH_X1 port map( G => n13148
                           , D => n13238, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_9_21_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_9_19_inst : DLH_X1 port map( G => n17714
                           , D => n13232, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_9_19_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_9_17_inst : DLH_X1 port map( G => n13148
                           , D => n13226, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_9_17_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_9_15_inst : DLH_X1 port map( G => n17714
                           , D => n13220, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_9_15_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_9_13_inst : DLH_X1 port map( G => n13148
                           , D => n13214, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_9_13_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_9_0_inst : DLH_X1 port map( G => n17714,
                           D => n13175, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_9_0_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_9_8_inst : DLH_X1 port map( G => n17714,
                           D => n13199, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_9_8_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_9_14_inst : DLH_X1 port map( G => n13148
                           , D => n13217, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_9_14_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_9_16_inst : DLH_X1 port map( G => n17714
                           , D => n13223, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_9_16_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_9_18_inst : DLH_X1 port map( G => n17714
                           , D => n13229, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_9_18_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_9_20_inst : DLH_X1 port map( G => n13148
                           , D => n13235, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_9_20_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_9_22_inst : DLH_X1 port map( G => n13148
                           , D => n13241, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_9_22_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_9_24_inst : DLH_X1 port map( G => n13148
                           , D => n13247, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_9_24_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_9_26_inst : DLH_X1 port map( G => n13148
                           , D => n13253, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_9_26_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_9_28_inst : DLH_X1 port map( G => n13148
                           , D => n13259, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_9_28_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_9_30_inst : DLH_X1 port map( G => n17714
                           , D => n13265, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_9_30_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_10_31_inst : DLH_X1 port map( G => 
                           n13145, D => n13268, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_10_31_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_10_29_inst : DLH_X1 port map( G => 
                           n17715, D => n13262, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_10_29_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_10_27_inst : DLH_X1 port map( G => 
                           n13145, D => n13256, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_10_27_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_10_25_inst : DLH_X1 port map( G => 
                           n17715, D => n13250, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_10_25_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_10_23_inst : DLH_X1 port map( G => 
                           n17715, D => n13244, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_10_23_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_10_21_inst : DLH_X1 port map( G => 
                           n13145, D => n13238, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_10_21_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_10_19_inst : DLH_X1 port map( G => 
                           n17715, D => n13232, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_10_19_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_10_17_inst : DLH_X1 port map( G => 
                           n13145, D => n13226, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_10_17_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_10_15_inst : DLH_X1 port map( G => 
                           n17715, D => n13220, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_10_15_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_10_13_inst : DLH_X1 port map( G => 
                           n13145, D => n13214, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_10_13_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_10_0_inst : DLH_X1 port map( G => n17715
                           , D => n13175, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_10_0_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_10_8_inst : DLH_X1 port map( G => n17715
                           , D => n13199, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_10_8_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_10_14_inst : DLH_X1 port map( G => 
                           n13145, D => n13217, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_10_14_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_10_16_inst : DLH_X1 port map( G => 
                           n17715, D => n13223, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_10_16_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_10_18_inst : DLH_X1 port map( G => 
                           n17715, D => n13229, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_10_18_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_10_20_inst : DLH_X1 port map( G => 
                           n13145, D => n13235, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_10_20_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_10_22_inst : DLH_X1 port map( G => 
                           n13145, D => n13241, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_10_22_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_10_24_inst : DLH_X1 port map( G => 
                           n13145, D => n13247, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_10_24_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_10_26_inst : DLH_X1 port map( G => 
                           n13145, D => n13253, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_10_26_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_10_28_inst : DLH_X1 port map( G => 
                           n13145, D => n13259, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_10_28_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_10_30_inst : DLH_X1 port map( G => 
                           n17715, D => n13265, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_10_30_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_11_31_inst : DLH_X1 port map( G => 
                           n13142, D => n13268, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_11_31_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_11_29_inst : DLH_X1 port map( G => 
                           n17716, D => n13262, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_11_29_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_11_27_inst : DLH_X1 port map( G => 
                           n13142, D => n13256, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_11_27_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_11_25_inst : DLH_X1 port map( G => 
                           n17716, D => n13250, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_11_25_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_11_23_inst : DLH_X1 port map( G => 
                           n17716, D => n13244, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_11_23_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_11_21_inst : DLH_X1 port map( G => 
                           n13142, D => n13238, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_11_21_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_11_19_inst : DLH_X1 port map( G => 
                           n17716, D => n13232, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_11_19_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_11_17_inst : DLH_X1 port map( G => 
                           n13142, D => n13226, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_11_17_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_11_15_inst : DLH_X1 port map( G => 
                           n17716, D => n13220, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_11_15_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_11_13_inst : DLH_X1 port map( G => 
                           n13142, D => n13214, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_11_13_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_11_0_inst : DLH_X1 port map( G => n17716
                           , D => n13175, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_11_0_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_11_8_inst : DLH_X1 port map( G => n17716
                           , D => n13199, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_11_8_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_11_14_inst : DLH_X1 port map( G => 
                           n13142, D => n13217, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_11_14_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_11_16_inst : DLH_X1 port map( G => 
                           n17716, D => n13223, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_11_16_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_11_18_inst : DLH_X1 port map( G => 
                           n17716, D => n13229, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_11_18_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_11_20_inst : DLH_X1 port map( G => 
                           n13142, D => n13235, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_11_20_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_11_22_inst : DLH_X1 port map( G => 
                           n13142, D => n13241, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_11_22_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_11_24_inst : DLH_X1 port map( G => 
                           n13142, D => n13247, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_11_24_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_11_26_inst : DLH_X1 port map( G => 
                           n13142, D => n13253, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_11_26_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_11_28_inst : DLH_X1 port map( G => 
                           n13142, D => n13259, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_11_28_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_11_30_inst : DLH_X1 port map( G => 
                           n17716, D => n13265, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_11_30_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_12_31_inst : DLH_X1 port map( G => 
                           n13139, D => n13268, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_12_31_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_12_29_inst : DLH_X1 port map( G => 
                           n17717, D => n13262, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_12_29_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_12_27_inst : DLH_X1 port map( G => 
                           n13139, D => n13256, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_12_27_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_12_25_inst : DLH_X1 port map( G => 
                           n17717, D => n13250, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_12_25_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_12_23_inst : DLH_X1 port map( G => 
                           n17717, D => n13244, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_12_23_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_12_21_inst : DLH_X1 port map( G => 
                           n13139, D => n13238, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_12_21_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_12_19_inst : DLH_X1 port map( G => 
                           n17717, D => n13232, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_12_19_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_12_17_inst : DLH_X1 port map( G => 
                           n13139, D => n13226, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_12_17_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_12_15_inst : DLH_X1 port map( G => 
                           n17717, D => n13220, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_12_15_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_12_13_inst : DLH_X1 port map( G => 
                           n13139, D => n13214, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_12_13_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_12_0_inst : DLH_X1 port map( G => n17717
                           , D => n13175, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_12_0_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_12_8_inst : DLH_X1 port map( G => n17717
                           , D => n13199, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_12_8_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_12_14_inst : DLH_X1 port map( G => 
                           n13139, D => n13217, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_12_14_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_12_16_inst : DLH_X1 port map( G => 
                           n17717, D => n13223, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_12_16_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_12_18_inst : DLH_X1 port map( G => 
                           n17717, D => n13229, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_12_18_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_12_20_inst : DLH_X1 port map( G => 
                           n13139, D => n13235, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_12_20_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_12_22_inst : DLH_X1 port map( G => 
                           n13139, D => n13241, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_12_22_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_12_24_inst : DLH_X1 port map( G => 
                           n13139, D => n13247, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_12_24_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_12_26_inst : DLH_X1 port map( G => 
                           n13139, D => n13253, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_12_26_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_12_28_inst : DLH_X1 port map( G => 
                           n13139, D => n13259, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_12_28_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_12_30_inst : DLH_X1 port map( G => 
                           n17717, D => n13265, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_12_30_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_13_31_inst : DLH_X1 port map( G => 
                           n13136, D => n13268, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_13_31_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_13_29_inst : DLH_X1 port map( G => 
                           n17718, D => n13262, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_13_29_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_13_27_inst : DLH_X1 port map( G => 
                           n13136, D => n13256, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_13_27_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_13_25_inst : DLH_X1 port map( G => 
                           n17718, D => n13250, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_13_25_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_13_23_inst : DLH_X1 port map( G => 
                           n17718, D => n13244, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_13_23_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_13_21_inst : DLH_X1 port map( G => 
                           n13136, D => n13238, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_13_21_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_13_19_inst : DLH_X1 port map( G => 
                           n17718, D => n13232, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_13_19_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_13_17_inst : DLH_X1 port map( G => 
                           n13136, D => n13226, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_13_17_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_13_15_inst : DLH_X1 port map( G => 
                           n17718, D => n13220, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_13_15_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_13_13_inst : DLH_X1 port map( G => 
                           n13136, D => n13214, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_13_13_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_13_0_inst : DLH_X1 port map( G => n17718
                           , D => n13175, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_13_0_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_13_8_inst : DLH_X1 port map( G => n17718
                           , D => n13199, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_13_8_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_13_14_inst : DLH_X1 port map( G => 
                           n13136, D => n13217, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_13_14_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_13_16_inst : DLH_X1 port map( G => 
                           n17718, D => n13223, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_13_16_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_13_18_inst : DLH_X1 port map( G => 
                           n17718, D => n13229, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_13_18_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_13_20_inst : DLH_X1 port map( G => 
                           n13136, D => n13235, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_13_20_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_13_22_inst : DLH_X1 port map( G => 
                           n13136, D => n13241, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_13_22_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_13_24_inst : DLH_X1 port map( G => 
                           n13136, D => n13247, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_13_24_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_13_26_inst : DLH_X1 port map( G => 
                           n13136, D => n13253, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_13_26_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_13_28_inst : DLH_X1 port map( G => 
                           n13136, D => n13259, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_13_28_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_13_30_inst : DLH_X1 port map( G => 
                           n17718, D => n13265, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_13_30_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_14_31_inst : DLH_X1 port map( G => 
                           n13133, D => n13268, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_14_31_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_14_29_inst : DLH_X1 port map( G => 
                           n17719, D => n13262, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_14_29_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_14_27_inst : DLH_X1 port map( G => 
                           n13133, D => n13256, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_14_27_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_14_25_inst : DLH_X1 port map( G => 
                           n17719, D => n13250, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_14_25_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_14_23_inst : DLH_X1 port map( G => 
                           n17719, D => n13244, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_14_23_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_14_21_inst : DLH_X1 port map( G => 
                           n13133, D => n13238, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_14_21_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_14_19_inst : DLH_X1 port map( G => 
                           n17719, D => n13232, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_14_19_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_14_17_inst : DLH_X1 port map( G => 
                           n13133, D => n13226, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_14_17_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_14_15_inst : DLH_X1 port map( G => 
                           n17719, D => n13220, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_14_15_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_14_13_inst : DLH_X1 port map( G => 
                           n13133, D => n13214, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_14_13_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_14_0_inst : DLH_X1 port map( G => n17719
                           , D => n13175, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_14_0_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_14_8_inst : DLH_X1 port map( G => n17719
                           , D => n13199, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_14_8_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_14_14_inst : DLH_X1 port map( G => 
                           n13133, D => n13217, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_14_14_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_14_16_inst : DLH_X1 port map( G => 
                           n17719, D => n13223, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_14_16_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_14_18_inst : DLH_X1 port map( G => 
                           n17719, D => n13229, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_14_18_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_14_20_inst : DLH_X1 port map( G => 
                           n13133, D => n13235, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_14_20_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_14_22_inst : DLH_X1 port map( G => 
                           n13133, D => n13241, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_14_22_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_14_24_inst : DLH_X1 port map( G => 
                           n13133, D => n13247, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_14_24_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_14_26_inst : DLH_X1 port map( G => 
                           n13133, D => n13253, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_14_26_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_14_28_inst : DLH_X1 port map( G => 
                           n13133, D => n13259, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_14_28_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_14_30_inst : DLH_X1 port map( G => 
                           n17719, D => n13265, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_14_30_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_15_31_inst : DLH_X1 port map( G => 
                           n13130, D => n13268, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_15_31_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_15_29_inst : DLH_X1 port map( G => 
                           n17720, D => n13262, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_15_29_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_15_27_inst : DLH_X1 port map( G => 
                           n13130, D => n13256, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_15_27_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_15_25_inst : DLH_X1 port map( G => 
                           n17720, D => n13250, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_15_25_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_15_23_inst : DLH_X1 port map( G => 
                           n17720, D => n13244, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_15_23_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_15_21_inst : DLH_X1 port map( G => 
                           n13130, D => n13238, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_15_21_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_15_19_inst : DLH_X1 port map( G => 
                           n17720, D => n13232, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_15_19_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_15_17_inst : DLH_X1 port map( G => 
                           n13130, D => n13226, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_15_17_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_15_15_inst : DLH_X1 port map( G => 
                           n17720, D => n13220, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_15_15_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_15_13_inst : DLH_X1 port map( G => 
                           n13130, D => n13214, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_15_13_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_15_0_inst : DLH_X1 port map( G => n17720
                           , D => n13175, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_15_0_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_15_8_inst : DLH_X1 port map( G => n17720
                           , D => n13199, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_15_8_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_15_14_inst : DLH_X1 port map( G => 
                           n13130, D => n13217, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_15_14_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_15_16_inst : DLH_X1 port map( G => 
                           n17720, D => n13223, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_15_16_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_15_18_inst : DLH_X1 port map( G => 
                           n17720, D => n13229, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_15_18_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_15_20_inst : DLH_X1 port map( G => 
                           n13130, D => n13235, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_15_20_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_15_22_inst : DLH_X1 port map( G => 
                           n13130, D => n13241, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_15_22_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_15_24_inst : DLH_X1 port map( G => 
                           n13130, D => n13247, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_15_24_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_15_26_inst : DLH_X1 port map( G => 
                           n13130, D => n13253, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_15_26_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_15_28_inst : DLH_X1 port map( G => 
                           n13130, D => n13259, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_15_28_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_15_30_inst : DLH_X1 port map( G => 
                           n17720, D => n13265, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_15_30_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_16_31_inst : DLH_X1 port map( G => 
                           n13127, D => n13268, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_16_31_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_16_29_inst : DLH_X1 port map( G => 
                           n17721, D => n13262, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_16_29_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_16_27_inst : DLH_X1 port map( G => 
                           n13127, D => n13256, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_16_27_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_16_25_inst : DLH_X1 port map( G => 
                           n17721, D => n13250, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_16_25_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_16_23_inst : DLH_X1 port map( G => 
                           n17721, D => n13244, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_16_23_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_16_21_inst : DLH_X1 port map( G => 
                           n13127, D => n13238, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_16_21_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_16_19_inst : DLH_X1 port map( G => 
                           n17721, D => n13232, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_16_19_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_16_17_inst : DLH_X1 port map( G => 
                           n13127, D => n13226, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_16_17_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_16_15_inst : DLH_X1 port map( G => 
                           n17721, D => n13220, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_16_15_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_16_13_inst : DLH_X1 port map( G => 
                           n13127, D => n13214, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_16_13_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_16_0_inst : DLH_X1 port map( G => n17721
                           , D => n13175, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_16_0_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_16_8_inst : DLH_X1 port map( G => n17721
                           , D => n13199, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_16_8_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_16_14_inst : DLH_X1 port map( G => 
                           n13127, D => n13217, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_16_14_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_16_16_inst : DLH_X1 port map( G => 
                           n17721, D => n13223, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_16_16_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_16_18_inst : DLH_X1 port map( G => 
                           n17721, D => n13229, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_16_18_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_16_20_inst : DLH_X1 port map( G => 
                           n13127, D => n13235, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_16_20_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_16_22_inst : DLH_X1 port map( G => 
                           n13127, D => n13241, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_16_22_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_16_24_inst : DLH_X1 port map( G => 
                           n13127, D => n13247, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_16_24_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_16_26_inst : DLH_X1 port map( G => 
                           n13127, D => n13253, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_16_26_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_16_28_inst : DLH_X1 port map( G => 
                           n13127, D => n13259, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_16_28_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_16_30_inst : DLH_X1 port map( G => 
                           n17721, D => n13265, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_16_30_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_17_31_inst : DLH_X1 port map( G => 
                           n13124, D => n13268, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_17_31_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_17_29_inst : DLH_X1 port map( G => 
                           n17722, D => n13262, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_17_29_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_17_27_inst : DLH_X1 port map( G => 
                           n13124, D => n13256, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_17_27_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_17_25_inst : DLH_X1 port map( G => 
                           n17722, D => n13250, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_17_25_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_17_23_inst : DLH_X1 port map( G => 
                           n17722, D => n13244, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_17_23_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_17_21_inst : DLH_X1 port map( G => 
                           n13124, D => n13238, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_17_21_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_17_19_inst : DLH_X1 port map( G => 
                           n17722, D => n13232, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_17_19_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_17_17_inst : DLH_X1 port map( G => 
                           n13124, D => n13226, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_17_17_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_17_15_inst : DLH_X1 port map( G => 
                           n17722, D => n13220, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_17_15_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_17_13_inst : DLH_X1 port map( G => 
                           n13124, D => n13214, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_17_13_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_17_0_inst : DLH_X1 port map( G => n17722
                           , D => n13175, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_17_0_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_17_8_inst : DLH_X1 port map( G => n17722
                           , D => n13199, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_17_8_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_17_14_inst : DLH_X1 port map( G => 
                           n13124, D => n13217, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_17_14_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_17_16_inst : DLH_X1 port map( G => 
                           n17722, D => n13223, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_17_16_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_17_18_inst : DLH_X1 port map( G => 
                           n17722, D => n13229, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_17_18_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_17_20_inst : DLH_X1 port map( G => 
                           n13124, D => n13235, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_17_20_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_17_22_inst : DLH_X1 port map( G => 
                           n13124, D => n13241, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_17_22_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_17_24_inst : DLH_X1 port map( G => 
                           n13124, D => n13247, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_17_24_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_17_26_inst : DLH_X1 port map( G => 
                           n13124, D => n13253, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_17_26_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_17_28_inst : DLH_X1 port map( G => 
                           n13124, D => n13259, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_17_28_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_17_30_inst : DLH_X1 port map( G => 
                           n17722, D => n13265, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_17_30_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_18_31_inst : DLH_X1 port map( G => 
                           n13121, D => n13268, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_18_31_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_18_29_inst : DLH_X1 port map( G => 
                           n17723, D => n13262, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_18_29_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_18_27_inst : DLH_X1 port map( G => 
                           n13121, D => n13256, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_18_27_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_18_25_inst : DLH_X1 port map( G => 
                           n17723, D => n13250, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_18_25_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_18_23_inst : DLH_X1 port map( G => 
                           n17723, D => n13244, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_18_23_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_18_21_inst : DLH_X1 port map( G => 
                           n13121, D => n13238, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_18_21_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_18_19_inst : DLH_X1 port map( G => 
                           n17723, D => n13232, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_18_19_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_18_17_inst : DLH_X1 port map( G => 
                           n13121, D => n13226, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_18_17_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_18_15_inst : DLH_X1 port map( G => 
                           n17723, D => n13220, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_18_15_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_18_13_inst : DLH_X1 port map( G => 
                           n13121, D => n13214, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_18_13_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_18_0_inst : DLH_X1 port map( G => n17723
                           , D => n13175, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_18_0_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_18_8_inst : DLH_X1 port map( G => n17723
                           , D => n13199, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_18_8_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_18_14_inst : DLH_X1 port map( G => 
                           n13121, D => n13217, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_18_14_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_18_16_inst : DLH_X1 port map( G => 
                           n17723, D => n13223, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_18_16_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_18_18_inst : DLH_X1 port map( G => 
                           n17723, D => n13229, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_18_18_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_18_20_inst : DLH_X1 port map( G => 
                           n13121, D => n13235, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_18_20_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_18_22_inst : DLH_X1 port map( G => 
                           n13121, D => n13241, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_18_22_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_18_24_inst : DLH_X1 port map( G => 
                           n13121, D => n13247, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_18_24_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_18_26_inst : DLH_X1 port map( G => 
                           n13121, D => n13253, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_18_26_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_18_28_inst : DLH_X1 port map( G => 
                           n13121, D => n13259, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_18_28_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_18_30_inst : DLH_X1 port map( G => 
                           n17723, D => n13265, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_18_30_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_19_31_inst : DLH_X1 port map( G => 
                           n13118, D => n13268, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_19_31_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_19_29_inst : DLH_X1 port map( G => 
                           n17724, D => n13262, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_19_29_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_19_27_inst : DLH_X1 port map( G => 
                           n13118, D => n13256, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_19_27_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_19_25_inst : DLH_X1 port map( G => 
                           n17724, D => n13250, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_19_25_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_19_23_inst : DLH_X1 port map( G => 
                           n17724, D => n13244, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_19_23_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_19_21_inst : DLH_X1 port map( G => 
                           n13118, D => n13238, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_19_21_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_19_19_inst : DLH_X1 port map( G => 
                           n17724, D => n13232, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_19_19_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_19_17_inst : DLH_X1 port map( G => 
                           n13118, D => n13226, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_19_17_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_19_15_inst : DLH_X1 port map( G => 
                           n17724, D => n13220, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_19_15_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_19_13_inst : DLH_X1 port map( G => 
                           n13118, D => n13214, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_19_13_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_19_0_inst : DLH_X1 port map( G => n17724
                           , D => n13175, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_19_0_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_19_8_inst : DLH_X1 port map( G => n17724
                           , D => n13199, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_19_8_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_19_14_inst : DLH_X1 port map( G => 
                           n13118, D => n13217, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_19_14_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_19_16_inst : DLH_X1 port map( G => 
                           n17724, D => n13223, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_19_16_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_19_18_inst : DLH_X1 port map( G => 
                           n17724, D => n13229, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_19_18_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_19_20_inst : DLH_X1 port map( G => 
                           n13118, D => n13235, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_19_20_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_19_22_inst : DLH_X1 port map( G => 
                           n13118, D => n13241, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_19_22_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_19_24_inst : DLH_X1 port map( G => 
                           n13118, D => n13247, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_19_24_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_19_26_inst : DLH_X1 port map( G => 
                           n13118, D => n13253, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_19_26_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_19_28_inst : DLH_X1 port map( G => 
                           n13118, D => n13259, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_19_28_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_19_30_inst : DLH_X1 port map( G => 
                           n17724, D => n13265, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_19_30_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_20_31_inst : DLH_X1 port map( G => 
                           n13115, D => n13268, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_20_31_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_20_29_inst : DLH_X1 port map( G => 
                           n17725, D => n13262, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_20_29_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_20_27_inst : DLH_X1 port map( G => 
                           n13115, D => n13256, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_20_27_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_20_25_inst : DLH_X1 port map( G => 
                           n17725, D => n13250, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_20_25_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_20_23_inst : DLH_X1 port map( G => 
                           n17725, D => n13244, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_20_23_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_20_21_inst : DLH_X1 port map( G => 
                           n13115, D => n13238, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_20_21_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_20_19_inst : DLH_X1 port map( G => 
                           n17725, D => n13232, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_20_19_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_20_17_inst : DLH_X1 port map( G => 
                           n13115, D => n13226, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_20_17_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_20_15_inst : DLH_X1 port map( G => 
                           n17725, D => n13220, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_20_15_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_20_13_inst : DLH_X1 port map( G => 
                           n13115, D => n13214, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_20_13_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_20_0_inst : DLH_X1 port map( G => n17725
                           , D => n13175, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_20_0_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_20_8_inst : DLH_X1 port map( G => n17725
                           , D => n13199, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_20_8_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_20_14_inst : DLH_X1 port map( G => 
                           n13115, D => n13217, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_20_14_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_20_16_inst : DLH_X1 port map( G => 
                           n17725, D => n13223, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_20_16_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_20_18_inst : DLH_X1 port map( G => 
                           n17725, D => n13229, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_20_18_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_20_20_inst : DLH_X1 port map( G => 
                           n13115, D => n13235, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_20_20_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_20_22_inst : DLH_X1 port map( G => 
                           n13115, D => n13241, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_20_22_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_20_24_inst : DLH_X1 port map( G => 
                           n13115, D => n13247, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_20_24_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_20_26_inst : DLH_X1 port map( G => 
                           n13115, D => n13253, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_20_26_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_20_28_inst : DLH_X1 port map( G => 
                           n13115, D => n13259, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_20_28_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_20_30_inst : DLH_X1 port map( G => 
                           n17725, D => n13265, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_20_30_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_21_31_inst : DLH_X1 port map( G => 
                           n13112, D => n13268, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_21_31_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_21_29_inst : DLH_X1 port map( G => 
                           n17726, D => n13262, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_21_29_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_21_27_inst : DLH_X1 port map( G => 
                           n13112, D => n13256, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_21_27_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_21_25_inst : DLH_X1 port map( G => 
                           n17726, D => n13250, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_21_25_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_21_23_inst : DLH_X1 port map( G => 
                           n17726, D => n13244, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_21_23_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_21_21_inst : DLH_X1 port map( G => 
                           n13112, D => n13238, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_21_21_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_21_19_inst : DLH_X1 port map( G => 
                           n17726, D => n13232, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_21_19_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_21_17_inst : DLH_X1 port map( G => 
                           n13112, D => n13226, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_21_17_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_21_15_inst : DLH_X1 port map( G => 
                           n17726, D => n13220, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_21_15_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_21_13_inst : DLH_X1 port map( G => 
                           n13112, D => n13214, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_21_13_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_21_0_inst : DLH_X1 port map( G => n17726
                           , D => n13175, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_21_0_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_21_8_inst : DLH_X1 port map( G => n17726
                           , D => n13199, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_21_8_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_21_14_inst : DLH_X1 port map( G => 
                           n13112, D => n13217, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_21_14_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_21_16_inst : DLH_X1 port map( G => 
                           n17726, D => n13223, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_21_16_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_21_18_inst : DLH_X1 port map( G => 
                           n17726, D => n13229, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_21_18_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_21_20_inst : DLH_X1 port map( G => 
                           n13112, D => n13235, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_21_20_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_21_22_inst : DLH_X1 port map( G => 
                           n13112, D => n13241, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_21_22_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_21_24_inst : DLH_X1 port map( G => 
                           n13112, D => n13247, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_21_24_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_21_26_inst : DLH_X1 port map( G => 
                           n13112, D => n13253, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_21_26_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_21_28_inst : DLH_X1 port map( G => 
                           n13112, D => n13259, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_21_28_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_21_30_inst : DLH_X1 port map( G => 
                           n17726, D => n13265, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_21_30_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_22_31_inst : DLH_X1 port map( G => 
                           n13109, D => n13268, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_22_31_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_22_29_inst : DLH_X1 port map( G => 
                           n17727, D => n13262, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_22_29_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_22_27_inst : DLH_X1 port map( G => 
                           n13109, D => n13256, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_22_27_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_22_25_inst : DLH_X1 port map( G => 
                           n17727, D => n13250, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_22_25_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_22_23_inst : DLH_X1 port map( G => 
                           n17727, D => n13244, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_22_23_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_22_21_inst : DLH_X1 port map( G => 
                           n13109, D => n13238, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_22_21_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_22_19_inst : DLH_X1 port map( G => 
                           n17727, D => n13232, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_22_19_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_22_17_inst : DLH_X1 port map( G => 
                           n13109, D => n13226, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_22_17_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_22_15_inst : DLH_X1 port map( G => 
                           n17727, D => n13220, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_22_15_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_22_13_inst : DLH_X1 port map( G => 
                           n13109, D => n13214, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_22_13_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_22_0_inst : DLH_X1 port map( G => n17727
                           , D => n13175, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_22_0_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_22_8_inst : DLH_X1 port map( G => n17727
                           , D => n13199, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_22_8_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_22_14_inst : DLH_X1 port map( G => 
                           n13109, D => n13217, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_22_14_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_22_16_inst : DLH_X1 port map( G => 
                           n17727, D => n13223, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_22_16_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_22_18_inst : DLH_X1 port map( G => 
                           n17727, D => n13229, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_22_18_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_22_20_inst : DLH_X1 port map( G => 
                           n13109, D => n13235, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_22_20_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_22_22_inst : DLH_X1 port map( G => 
                           n13109, D => n13241, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_22_22_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_22_24_inst : DLH_X1 port map( G => 
                           n13109, D => n13247, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_22_24_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_22_26_inst : DLH_X1 port map( G => 
                           n13109, D => n13253, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_22_26_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_22_28_inst : DLH_X1 port map( G => 
                           n13109, D => n13259, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_22_28_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_22_30_inst : DLH_X1 port map( G => 
                           n17727, D => n13265, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_22_30_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_23_31_inst : DLH_X1 port map( G => 
                           n13106, D => n13268, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_23_31_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_23_29_inst : DLH_X1 port map( G => 
                           n17728, D => n13262, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_23_29_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_23_27_inst : DLH_X1 port map( G => 
                           n13106, D => n13256, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_23_27_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_23_25_inst : DLH_X1 port map( G => 
                           n17728, D => n13250, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_23_25_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_23_23_inst : DLH_X1 port map( G => 
                           n17728, D => n13244, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_23_23_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_23_21_inst : DLH_X1 port map( G => 
                           n13106, D => n13238, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_23_21_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_23_19_inst : DLH_X1 port map( G => 
                           n17728, D => n13232, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_23_19_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_23_17_inst : DLH_X1 port map( G => 
                           n13106, D => n13226, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_23_17_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_23_15_inst : DLH_X1 port map( G => 
                           n17728, D => n13220, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_23_15_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_23_13_inst : DLH_X1 port map( G => 
                           n13106, D => n13214, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_23_13_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_23_0_inst : DLH_X1 port map( G => n17728
                           , D => n13175, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_23_0_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_23_8_inst : DLH_X1 port map( G => n17728
                           , D => n13199, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_23_8_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_23_14_inst : DLH_X1 port map( G => 
                           n13106, D => n13217, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_23_14_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_23_16_inst : DLH_X1 port map( G => 
                           n17728, D => n13223, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_23_16_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_23_18_inst : DLH_X1 port map( G => 
                           n17728, D => n13229, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_23_18_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_23_20_inst : DLH_X1 port map( G => 
                           n13106, D => n13235, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_23_20_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_23_22_inst : DLH_X1 port map( G => 
                           n13106, D => n13241, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_23_22_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_23_24_inst : DLH_X1 port map( G => 
                           n13106, D => n13247, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_23_24_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_23_26_inst : DLH_X1 port map( G => 
                           n13106, D => n13253, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_23_26_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_23_28_inst : DLH_X1 port map( G => 
                           n13106, D => n13259, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_23_28_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_23_30_inst : DLH_X1 port map( G => 
                           n17728, D => n13265, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_23_30_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_24_31_inst : DLH_X1 port map( G => 
                           n13103, D => n13268, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_24_31_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_24_29_inst : DLH_X1 port map( G => 
                           n17729, D => n13262, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_24_29_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_24_27_inst : DLH_X1 port map( G => 
                           n13103, D => n13256, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_24_27_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_24_25_inst : DLH_X1 port map( G => 
                           n17729, D => n13250, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_24_25_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_24_23_inst : DLH_X1 port map( G => 
                           n17729, D => n13244, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_24_23_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_24_21_inst : DLH_X1 port map( G => 
                           n13103, D => n13238, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_24_21_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_24_19_inst : DLH_X1 port map( G => 
                           n17729, D => n13232, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_24_19_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_24_17_inst : DLH_X1 port map( G => 
                           n13103, D => n13226, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_24_17_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_24_15_inst : DLH_X1 port map( G => 
                           n17729, D => n13220, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_24_15_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_24_13_inst : DLH_X1 port map( G => 
                           n13103, D => n13214, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_24_13_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_24_0_inst : DLH_X1 port map( G => n17729
                           , D => n13175, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_24_0_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_24_8_inst : DLH_X1 port map( G => n17729
                           , D => n13199, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_24_8_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_24_14_inst : DLH_X1 port map( G => 
                           n13103, D => n13217, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_24_14_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_24_16_inst : DLH_X1 port map( G => 
                           n17729, D => n13223, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_24_16_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_24_18_inst : DLH_X1 port map( G => 
                           n17729, D => n13229, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_24_18_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_24_20_inst : DLH_X1 port map( G => 
                           n13103, D => n13235, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_24_20_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_24_22_inst : DLH_X1 port map( G => 
                           n13103, D => n13241, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_24_22_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_24_24_inst : DLH_X1 port map( G => 
                           n13103, D => n13247, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_24_24_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_24_26_inst : DLH_X1 port map( G => 
                           n13103, D => n13253, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_24_26_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_24_28_inst : DLH_X1 port map( G => 
                           n13103, D => n13259, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_24_28_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_24_30_inst : DLH_X1 port map( G => 
                           n17729, D => n13265, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_24_30_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_25_31_inst : DLH_X1 port map( G => 
                           n13100, D => n13268, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_25_31_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_25_29_inst : DLH_X1 port map( G => 
                           n17730, D => n13262, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_25_29_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_25_27_inst : DLH_X1 port map( G => 
                           n13100, D => n13256, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_25_27_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_25_25_inst : DLH_X1 port map( G => 
                           n17730, D => n13250, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_25_25_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_25_23_inst : DLH_X1 port map( G => 
                           n17730, D => n13244, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_25_23_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_25_21_inst : DLH_X1 port map( G => 
                           n13100, D => n13238, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_25_21_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_25_19_inst : DLH_X1 port map( G => 
                           n17730, D => n13232, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_25_19_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_25_17_inst : DLH_X1 port map( G => 
                           n13100, D => n13226, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_25_17_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_25_15_inst : DLH_X1 port map( G => 
                           n17730, D => n13220, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_25_15_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_25_13_inst : DLH_X1 port map( G => 
                           n13100, D => n13214, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_25_13_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_25_0_inst : DLH_X1 port map( G => n17730
                           , D => n13175, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_25_0_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_25_8_inst : DLH_X1 port map( G => n17730
                           , D => n13199, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_25_8_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_25_14_inst : DLH_X1 port map( G => 
                           n13100, D => n13217, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_25_14_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_25_16_inst : DLH_X1 port map( G => 
                           n17730, D => n13223, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_25_16_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_25_18_inst : DLH_X1 port map( G => 
                           n17730, D => n13229, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_25_18_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_25_20_inst : DLH_X1 port map( G => 
                           n13100, D => n13235, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_25_20_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_25_22_inst : DLH_X1 port map( G => 
                           n13100, D => n13241, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_25_22_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_25_24_inst : DLH_X1 port map( G => 
                           n13100, D => n13247, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_25_24_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_25_26_inst : DLH_X1 port map( G => 
                           n13100, D => n13253, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_25_26_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_25_28_inst : DLH_X1 port map( G => 
                           n13100, D => n13259, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_25_28_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_25_30_inst : DLH_X1 port map( G => 
                           n17730, D => n13265, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_25_30_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_26_31_inst : DLH_X1 port map( G => 
                           n13097, D => n13268, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_26_31_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_26_29_inst : DLH_X1 port map( G => 
                           n17731, D => n13262, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_26_29_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_26_27_inst : DLH_X1 port map( G => 
                           n13097, D => n13256, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_26_27_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_26_25_inst : DLH_X1 port map( G => 
                           n17731, D => n13250, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_26_25_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_26_23_inst : DLH_X1 port map( G => 
                           n17731, D => n13244, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_26_23_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_26_21_inst : DLH_X1 port map( G => 
                           n13097, D => n13238, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_26_21_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_26_19_inst : DLH_X1 port map( G => 
                           n17731, D => n13232, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_26_19_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_26_17_inst : DLH_X1 port map( G => 
                           n13097, D => n13226, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_26_17_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_26_15_inst : DLH_X1 port map( G => 
                           n17731, D => n13220, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_26_15_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_26_13_inst : DLH_X1 port map( G => 
                           n13097, D => n13214, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_26_13_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_26_0_inst : DLH_X1 port map( G => n17731
                           , D => n13175, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_26_0_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_26_8_inst : DLH_X1 port map( G => n17731
                           , D => n13199, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_26_8_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_26_14_inst : DLH_X1 port map( G => 
                           n13097, D => n13217, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_26_14_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_26_16_inst : DLH_X1 port map( G => 
                           n17731, D => n13223, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_26_16_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_26_18_inst : DLH_X1 port map( G => 
                           n17731, D => n13229, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_26_18_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_26_20_inst : DLH_X1 port map( G => 
                           n13097, D => n13235, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_26_20_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_26_22_inst : DLH_X1 port map( G => 
                           n13097, D => n13241, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_26_22_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_26_24_inst : DLH_X1 port map( G => 
                           n13097, D => n13247, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_26_24_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_26_26_inst : DLH_X1 port map( G => 
                           n13097, D => n13253, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_26_26_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_26_28_inst : DLH_X1 port map( G => 
                           n13097, D => n13259, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_26_28_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_26_30_inst : DLH_X1 port map( G => 
                           n17731, D => n13265, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_26_30_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_27_31_inst : DLH_X1 port map( G => 
                           n13094, D => n13268, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_27_31_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_27_29_inst : DLH_X1 port map( G => 
                           n17732, D => n13262, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_27_29_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_27_27_inst : DLH_X1 port map( G => 
                           n13094, D => n13256, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_27_27_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_27_25_inst : DLH_X1 port map( G => 
                           n17732, D => n13250, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_27_25_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_27_23_inst : DLH_X1 port map( G => 
                           n17732, D => n13244, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_27_23_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_27_21_inst : DLH_X1 port map( G => 
                           n13094, D => n13238, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_27_21_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_27_19_inst : DLH_X1 port map( G => 
                           n17732, D => n13232, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_27_19_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_27_17_inst : DLH_X1 port map( G => 
                           n13094, D => n13226, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_27_17_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_27_15_inst : DLH_X1 port map( G => 
                           n17732, D => n13220, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_27_15_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_27_13_inst : DLH_X1 port map( G => 
                           n13094, D => n13214, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_27_13_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_27_0_inst : DLH_X1 port map( G => n17732
                           , D => n13175, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_27_0_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_27_8_inst : DLH_X1 port map( G => n17732
                           , D => n13199, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_27_8_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_27_14_inst : DLH_X1 port map( G => 
                           n13094, D => n13217, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_27_14_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_27_16_inst : DLH_X1 port map( G => 
                           n17732, D => n13223, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_27_16_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_27_18_inst : DLH_X1 port map( G => 
                           n17732, D => n13229, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_27_18_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_27_20_inst : DLH_X1 port map( G => 
                           n13094, D => n13235, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_27_20_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_27_22_inst : DLH_X1 port map( G => 
                           n13094, D => n13241, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_27_22_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_27_24_inst : DLH_X1 port map( G => 
                           n13094, D => n13247, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_27_24_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_27_26_inst : DLH_X1 port map( G => 
                           n13094, D => n13253, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_27_26_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_27_28_inst : DLH_X1 port map( G => 
                           n13094, D => n13259, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_27_28_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_27_30_inst : DLH_X1 port map( G => 
                           n17732, D => n13265, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_27_30_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_28_31_inst : DLH_X1 port map( G => 
                           n13091, D => n13268, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_28_31_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_28_29_inst : DLH_X1 port map( G => 
                           n17733, D => n13262, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_28_29_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_28_27_inst : DLH_X1 port map( G => 
                           n13091, D => n13256, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_28_27_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_28_25_inst : DLH_X1 port map( G => 
                           n17733, D => n13250, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_28_25_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_28_23_inst : DLH_X1 port map( G => 
                           n17733, D => n13244, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_28_23_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_28_21_inst : DLH_X1 port map( G => 
                           n13091, D => n13238, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_28_21_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_28_19_inst : DLH_X1 port map( G => 
                           n17733, D => n13232, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_28_19_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_28_17_inst : DLH_X1 port map( G => 
                           n13091, D => n13226, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_28_17_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_28_15_inst : DLH_X1 port map( G => 
                           n17733, D => n13220, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_28_15_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_28_13_inst : DLH_X1 port map( G => 
                           n13091, D => n13214, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_28_13_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_28_0_inst : DLH_X1 port map( G => n17733
                           , D => n13175, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_28_0_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_28_8_inst : DLH_X1 port map( G => n17733
                           , D => n13199, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_28_8_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_28_14_inst : DLH_X1 port map( G => 
                           n13091, D => n13217, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_28_14_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_28_16_inst : DLH_X1 port map( G => 
                           n17733, D => n13223, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_28_16_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_28_18_inst : DLH_X1 port map( G => 
                           n17733, D => n13229, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_28_18_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_28_20_inst : DLH_X1 port map( G => 
                           n13091, D => n13235, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_28_20_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_28_22_inst : DLH_X1 port map( G => 
                           n13091, D => n13241, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_28_22_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_28_24_inst : DLH_X1 port map( G => 
                           n13091, D => n13247, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_28_24_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_28_26_inst : DLH_X1 port map( G => 
                           n13091, D => n13253, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_28_26_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_28_28_inst : DLH_X1 port map( G => 
                           n13091, D => n13259, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_28_28_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_28_30_inst : DLH_X1 port map( G => 
                           n17733, D => n13265, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_28_30_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_29_31_inst : DLH_X1 port map( G => 
                           n13088, D => n13268, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_29_31_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_29_29_inst : DLH_X1 port map( G => 
                           n17734, D => n13262, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_29_29_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_29_27_inst : DLH_X1 port map( G => 
                           n13088, D => n13256, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_29_27_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_29_25_inst : DLH_X1 port map( G => 
                           n17734, D => n13250, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_29_25_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_29_23_inst : DLH_X1 port map( G => 
                           n17734, D => n13244, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_29_23_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_29_21_inst : DLH_X1 port map( G => 
                           n13088, D => n13238, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_29_21_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_29_19_inst : DLH_X1 port map( G => 
                           n17734, D => n13232, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_29_19_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_29_17_inst : DLH_X1 port map( G => 
                           n13088, D => n13226, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_29_17_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_29_15_inst : DLH_X1 port map( G => 
                           n17734, D => n13220, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_29_15_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_29_13_inst : DLH_X1 port map( G => 
                           n13088, D => n13214, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_29_13_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_29_0_inst : DLH_X1 port map( G => n17734
                           , D => n13175, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_29_0_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_29_8_inst : DLH_X1 port map( G => n17734
                           , D => n13199, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_29_8_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_29_14_inst : DLH_X1 port map( G => 
                           n13088, D => n13217, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_29_14_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_29_16_inst : DLH_X1 port map( G => 
                           n17734, D => n13223, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_29_16_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_29_18_inst : DLH_X1 port map( G => 
                           n17734, D => n13229, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_29_18_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_29_20_inst : DLH_X1 port map( G => 
                           n13088, D => n13235, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_29_20_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_29_22_inst : DLH_X1 port map( G => 
                           n13088, D => n13241, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_29_22_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_29_24_inst : DLH_X1 port map( G => 
                           n13088, D => n13247, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_29_24_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_29_26_inst : DLH_X1 port map( G => 
                           n13088, D => n13253, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_29_26_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_29_28_inst : DLH_X1 port map( G => 
                           n13088, D => n13259, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_29_28_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_29_30_inst : DLH_X1 port map( G => 
                           n17734, D => n13265, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_29_30_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_30_31_inst : DLH_X1 port map( G => 
                           n13085, D => n13268, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_30_31_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_30_29_inst : DLH_X1 port map( G => 
                           n17735, D => n13262, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_30_29_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_30_27_inst : DLH_X1 port map( G => 
                           n13085, D => n13256, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_30_27_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_30_25_inst : DLH_X1 port map( G => 
                           n17735, D => n13250, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_30_25_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_30_23_inst : DLH_X1 port map( G => 
                           n17735, D => n13244, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_30_23_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_30_21_inst : DLH_X1 port map( G => 
                           n13085, D => n13238, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_30_21_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_30_19_inst : DLH_X1 port map( G => 
                           n17735, D => n13232, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_30_19_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_30_17_inst : DLH_X1 port map( G => 
                           n13085, D => n13226, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_30_17_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_30_15_inst : DLH_X1 port map( G => 
                           n17735, D => n13220, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_30_15_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_30_13_inst : DLH_X1 port map( G => 
                           n13085, D => n13214, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_30_13_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_30_0_inst : DLH_X1 port map( G => n17735
                           , D => n13175, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_30_0_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_30_8_inst : DLH_X1 port map( G => n17735
                           , D => n13199, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_30_8_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_30_14_inst : DLH_X1 port map( G => 
                           n13085, D => n13217, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_30_14_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_30_16_inst : DLH_X1 port map( G => 
                           n17735, D => n13223, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_30_16_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_30_18_inst : DLH_X1 port map( G => 
                           n17735, D => n13229, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_30_18_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_30_20_inst : DLH_X1 port map( G => 
                           n13085, D => n13235, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_30_20_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_30_22_inst : DLH_X1 port map( G => 
                           n13085, D => n13241, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_30_22_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_30_24_inst : DLH_X1 port map( G => 
                           n13085, D => n13247, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_30_24_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_30_26_inst : DLH_X1 port map( G => 
                           n13085, D => n13253, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_30_26_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_30_28_inst : DLH_X1 port map( G => 
                           n13085, D => n13259, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_30_28_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_30_30_inst : DLH_X1 port map( G => 
                           n17735, D => n13265, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_30_30_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_31_31_inst : DLH_X1 port map( G => 
                           n13082, D => n13268, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_31_31_port);
   pipeline_IDEX_Stage_Reg2_out_IDEX_reg_31_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N165, CK => Clk, Q => n13886, QN
                           => n17526);
   pipeline_RegFile_DEC_WB_RegBank_reg_31_29_inst : DLH_X1 port map( G => 
                           n17736, D => n13262, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_31_29_port);
   pipeline_IDEX_Stage_Reg2_out_IDEX_reg_29_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N163, CK => Clk, Q => n13885, QN
                           => n17524);
   pipeline_RegFile_DEC_WB_RegBank_reg_31_27_inst : DLH_X1 port map( G => 
                           n13082, D => n13256, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_31_27_port);
   pipeline_IDEX_Stage_Reg2_out_IDEX_reg_27_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N161, CK => Clk, Q => n13884, QN
                           => n17522);
   pipeline_RegFile_DEC_WB_RegBank_reg_31_25_inst : DLH_X1 port map( G => 
                           n17736, D => n13250, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_31_25_port);
   pipeline_IDEX_Stage_Reg2_out_IDEX_reg_25_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N159, CK => Clk, Q => n13883, QN
                           => n17520);
   pipeline_RegFile_DEC_WB_RegBank_reg_31_23_inst : DLH_X1 port map( G => 
                           n17736, D => n13244, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_31_23_port);
   pipeline_IDEX_Stage_Reg2_out_IDEX_reg_23_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N157, CK => Clk, Q => n13882, QN
                           => n17518);
   pipeline_RegFile_DEC_WB_RegBank_reg_31_21_inst : DLH_X1 port map( G => 
                           n13082, D => n13238, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_31_21_port);
   pipeline_IDEX_Stage_Reg2_out_IDEX_reg_21_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N155, CK => Clk, Q => n13881, QN
                           => n17516);
   pipeline_RegFile_DEC_WB_RegBank_reg_31_19_inst : DLH_X1 port map( G => 
                           n17736, D => n13232, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_31_19_port);
   pipeline_IDEX_Stage_Reg2_out_IDEX_reg_19_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N153, CK => Clk, Q => n13880, QN
                           => n17514);
   pipeline_RegFile_DEC_WB_RegBank_reg_31_17_inst : DLH_X1 port map( G => 
                           n13082, D => n13226, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_31_17_port);
   pipeline_IDEX_Stage_Reg2_out_IDEX_reg_17_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N151, CK => Clk, Q => n13879, QN
                           => n17512);
   pipeline_RegFile_DEC_WB_RegBank_reg_31_15_inst : DLH_X1 port map( G => 
                           n17736, D => n13220, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_31_15_port);
   pipeline_IDEX_Stage_Reg2_out_IDEX_reg_15_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N149, CK => Clk, Q => n13878, QN
                           => n17510);
   pipeline_RegFile_DEC_WB_RegBank_reg_31_13_inst : DLH_X1 port map( G => 
                           n13082, D => n13214, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_31_13_port);
   pipeline_IDEX_Stage_Reg2_out_IDEX_reg_13_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N147, CK => Clk, Q => n13877, QN
                           => n17508);
   pipeline_RegFile_DEC_WB_RegBank_reg_31_0_inst : DLH_X1 port map( G => n17736
                           , D => n13175, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_31_0_port);
   pipeline_IDEX_Stage_Reg2_out_IDEX_reg_0_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N134, CK => Clk, Q => n13876, QN
                           => n17495);
   pipeline_RegFile_DEC_WB_RegBank_reg_31_8_inst : DLH_X1 port map( G => n17736
                           , D => n13199, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_31_8_port);
   pipeline_IDEX_Stage_Reg2_out_IDEX_reg_8_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N142, CK => Clk, Q => n13875, QN
                           => n17503);
   pipeline_RegFile_DEC_WB_RegBank_reg_31_14_inst : DLH_X1 port map( G => 
                           n13082, D => n13217, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_31_14_port);
   pipeline_IDEX_Stage_Reg2_out_IDEX_reg_14_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N148, CK => Clk, Q => n13874, QN
                           => n17509);
   pipeline_RegFile_DEC_WB_RegBank_reg_31_16_inst : DLH_X1 port map( G => 
                           n17736, D => n13223, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_31_16_port);
   pipeline_IDEX_Stage_Reg2_out_IDEX_reg_16_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N150, CK => Clk, Q => n13873, QN
                           => n17511);
   pipeline_RegFile_DEC_WB_RegBank_reg_31_18_inst : DLH_X1 port map( G => 
                           n17736, D => n13229, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_31_18_port);
   pipeline_IDEX_Stage_Reg2_out_IDEX_reg_18_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N152, CK => Clk, Q => n13872, QN
                           => n17513);
   pipeline_RegFile_DEC_WB_RegBank_reg_31_20_inst : DLH_X1 port map( G => 
                           n13082, D => n13235, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_31_20_port);
   pipeline_IDEX_Stage_Reg2_out_IDEX_reg_20_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N154, CK => Clk, Q => n13871, QN
                           => n17515);
   pipeline_RegFile_DEC_WB_RegBank_reg_31_22_inst : DLH_X1 port map( G => 
                           n13082, D => n13241, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_31_22_port);
   pipeline_IDEX_Stage_Reg2_out_IDEX_reg_22_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N156, CK => Clk, Q => n13870, QN
                           => n17517);
   pipeline_RegFile_DEC_WB_RegBank_reg_31_24_inst : DLH_X1 port map( G => 
                           n13082, D => n13247, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_31_24_port);
   pipeline_IDEX_Stage_Reg2_out_IDEX_reg_24_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N158, CK => Clk, Q => n13869, QN
                           => n17519);
   pipeline_RegFile_DEC_WB_RegBank_reg_31_26_inst : DLH_X1 port map( G => 
                           n13082, D => n13253, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_31_26_port);
   pipeline_IDEX_Stage_Reg2_out_IDEX_reg_26_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N160, CK => Clk, Q => n13868, QN
                           => n17521);
   pipeline_RegFile_DEC_WB_RegBank_reg_31_28_inst : DLH_X1 port map( G => 
                           n13082, D => n13259, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_31_28_port);
   pipeline_IDEX_Stage_Reg2_out_IDEX_reg_28_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N162, CK => Clk, Q => n13867, QN
                           => n17523);
   pipeline_RegFile_DEC_WB_RegBank_reg_31_30_inst : DLH_X1 port map( G => 
                           n17736, D => n13265, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_31_30_port);
   pipeline_IDEX_Stage_Reg2_out_IDEX_reg_30_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N164, CK => Clk, Q => n13866, QN
                           => n17525);
   pipeline_stageF_PC_reg_PC_out_reg_28_inst : DFFR_X1 port map( D => n3912, CK
                           => Clk, RN => n17705, Q => n13865, QN => n7675);
   pipeline_stageF_PC_reg_PC_out_reg_27_inst : DFFR_X1 port map( D => n3910, CK
                           => Clk, RN => n17703, Q => n13864, QN => n7674);
   pipeline_stageF_PC_reg_PC_out_reg_26_inst : DFFR_X1 port map( D => n3908, CK
                           => Clk, RN => n17702, Q => n13863, QN => n7673);
   pipeline_stageF_PC_reg_PC_out_reg_25_inst : DFFR_X1 port map( D => n3906, CK
                           => Clk, RN => n17705, Q => n13862, QN => n7672);
   pipeline_stageF_PC_reg_PC_out_reg_24_inst : DFFR_X1 port map( D => n3904, CK
                           => Clk, RN => n17705, Q => n13861, QN => n7671);
   pipeline_stageF_PC_reg_PC_out_reg_23_inst : DFFR_X1 port map( D => n3902, CK
                           => Clk, RN => n17705, Q => n13860, QN => n7670);
   pipeline_stageF_PC_reg_PC_out_reg_22_inst : DFFR_X1 port map( D => n3900, CK
                           => Clk, RN => n17703, Q => n13859, QN => n7669);
   pipeline_stageF_PC_reg_PC_out_reg_21_inst : DFFR_X1 port map( D => n3898, CK
                           => Clk, RN => n17705, Q => n13858, QN => n7668);
   pipeline_stageF_PC_reg_PC_out_reg_20_inst : DFFR_X1 port map( D => n3896, CK
                           => Clk, RN => n17705, Q => n13857, QN => n7667);
   pipeline_stageF_PC_reg_PC_out_reg_19_inst : DFFR_X1 port map( D => n3894, CK
                           => Clk, RN => n17704, Q => n13856, QN => n7666);
   pipeline_stageF_PC_reg_PC_out_reg_18_inst : DFFR_X1 port map( D => n3892, CK
                           => Clk, RN => n17705, Q => n13855, QN => n7665);
   pipeline_stageF_PC_reg_PC_out_reg_17_inst : DFFR_X1 port map( D => n3890, CK
                           => Clk, RN => n17705, Q => n13854, QN => n7664);
   pipeline_stageF_PC_reg_PC_out_reg_15_inst : DFFR_X1 port map( D => n3888, CK
                           => Clk, RN => n17705, Q => n13853, QN => n7663);
   pipeline_stageF_PC_reg_PC_out_reg_14_inst : DFFR_X1 port map( D => n3886, CK
                           => Clk, RN => n17705, Q => n13852, QN => n7662);
   pipeline_stageF_PC_reg_PC_out_reg_13_inst : DFFR_X1 port map( D => n3884, CK
                           => Clk, RN => n17701, Q => n13851, QN => n7661);
   pipeline_stageF_PC_reg_PC_out_reg_8_inst : DFFR_X1 port map( D => n3882, CK 
                           => Clk, RN => n17705, Q => n13850, QN => n7660);
   pipeline_stageF_PC_reg_PC_out_reg_0_inst : DFFR_X1 port map( D => n3880, CK 
                           => Clk, RN => n17704, Q => n13849, QN => n7659);
   DataMem_Mem_reg_0_1_inst : DLH_X1 port map( G => n13058, D => DataMem_N1651,
                           Q => DataMem_Mem_0_1_port);
   DataMem_Dataout_reg_1_inst : DLL_X1 port map( D => DataMem_N2164, GN => 
                           n17098, Q => DataMem_N2346);
   pipeline_MEMWB_Stage_Data_to_RF_reg_1_inst : DFF_X1 port map( D => 
                           pipeline_MEMWB_Stage_N12, CK => Clk, Q => 
                           pipeline_data_to_RF_from_WB_1_port, QN => n17321);
   pipeline_RegFile_DEC_WB_RegBank_reg_2_1_inst : DLH_X1 port map( G => n17707,
                           D => n13178, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_2_1_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_4_1_inst : DLH_X1 port map( G => n17709,
                           D => n13178, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_4_1_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_6_1_inst : DLH_X1 port map( G => n17711,
                           D => n13178, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_6_1_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_8_1_inst : DLH_X1 port map( G => n17713,
                           D => n13178, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_8_1_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_10_1_inst : DLH_X1 port map( G => n17715
                           , D => n13178, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_10_1_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_12_1_inst : DLH_X1 port map( G => n17717
                           , D => n13178, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_12_1_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_14_1_inst : DLH_X1 port map( G => n17719
                           , D => n13178, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_14_1_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_16_1_inst : DLH_X1 port map( G => n17721
                           , D => n13178, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_16_1_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_18_1_inst : DLH_X1 port map( G => n17723
                           , D => n13178, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_18_1_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_20_1_inst : DLH_X1 port map( G => n17725
                           , D => n13178, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_20_1_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_22_1_inst : DLH_X1 port map( G => n17727
                           , D => n13178, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_22_1_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_24_1_inst : DLH_X1 port map( G => n17729
                           , D => n13178, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_24_1_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_26_1_inst : DLH_X1 port map( G => n17731
                           , D => n13178, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_26_1_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_28_1_inst : DLH_X1 port map( G => n17733
                           , D => n13178, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_28_1_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_30_1_inst : DLH_X1 port map( G => n17735
                           , D => n13178, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_30_1_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_31_1_inst : DLH_X1 port map( G => n17736
                           , D => n13178, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_31_1_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_29_1_inst : DLH_X1 port map( G => n17734
                           , D => n13178, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_29_1_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_27_1_inst : DLH_X1 port map( G => n17732
                           , D => n13178, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_27_1_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_25_1_inst : DLH_X1 port map( G => n17730
                           , D => n13178, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_25_1_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_23_1_inst : DLH_X1 port map( G => n17728
                           , D => n13178, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_23_1_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_21_1_inst : DLH_X1 port map( G => n17726
                           , D => n13178, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_21_1_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_19_1_inst : DLH_X1 port map( G => n17724
                           , D => n13178, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_19_1_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_17_1_inst : DLH_X1 port map( G => n17722
                           , D => n13178, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_17_1_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_15_1_inst : DLH_X1 port map( G => n17720
                           , D => n13178, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_15_1_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_13_1_inst : DLH_X1 port map( G => n17718
                           , D => n13178, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_13_1_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_11_1_inst : DLH_X1 port map( G => n17716
                           , D => n13178, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_11_1_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_9_1_inst : DLH_X1 port map( G => n17714,
                           D => n13178, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_9_1_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_7_1_inst : DLH_X1 port map( G => n17712,
                           D => n13178, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_7_1_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_5_1_inst : DLH_X1 port map( G => n17710,
                           D => n13178, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_5_1_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_3_1_inst : DLH_X1 port map( G => n17708,
                           D => n13178, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_3_1_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_1_1_inst : DLH_X1 port map( G => n17706,
                           D => n13178, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_1_1_port);
   pipeline_IDEX_Stage_Reg2_out_IDEX_reg_1_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N135, CK => Clk, Q => n13848, QN
                           => n17496);
   pipeline_IDEX_Stage_Reg1_out_IDEX_reg_1_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N103, CK => Clk, Q => n13847, QN
                           => net214751);
   pipeline_MEMWB_Stage_Data_to_RF_reg_3_inst : DFF_X1 port map( D => 
                           pipeline_MEMWB_Stage_N14, CK => Clk, Q => 
                           pipeline_data_to_RF_from_WB_3_port, QN => n17306);
   pipeline_RegFile_DEC_WB_RegBank_reg_2_3_inst : DLH_X1 port map( G => n17707,
                           D => n13184, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_2_3_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_4_3_inst : DLH_X1 port map( G => n17709,
                           D => n13184, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_4_3_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_6_3_inst : DLH_X1 port map( G => n17711,
                           D => n13184, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_6_3_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_8_3_inst : DLH_X1 port map( G => n17713,
                           D => n13184, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_8_3_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_10_3_inst : DLH_X1 port map( G => n17715
                           , D => n13184, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_10_3_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_12_3_inst : DLH_X1 port map( G => n17717
                           , D => n13184, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_12_3_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_14_3_inst : DLH_X1 port map( G => n17719
                           , D => n13184, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_14_3_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_16_3_inst : DLH_X1 port map( G => n17721
                           , D => n13184, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_16_3_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_18_3_inst : DLH_X1 port map( G => n17723
                           , D => n13184, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_18_3_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_20_3_inst : DLH_X1 port map( G => n17725
                           , D => n13184, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_20_3_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_22_3_inst : DLH_X1 port map( G => n17727
                           , D => n13184, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_22_3_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_24_3_inst : DLH_X1 port map( G => n17729
                           , D => n13184, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_24_3_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_26_3_inst : DLH_X1 port map( G => n17731
                           , D => n13184, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_26_3_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_28_3_inst : DLH_X1 port map( G => n17733
                           , D => n13184, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_28_3_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_30_3_inst : DLH_X1 port map( G => n17735
                           , D => n13184, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_30_3_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_31_3_inst : DLH_X1 port map( G => n17736
                           , D => n13184, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_31_3_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_29_3_inst : DLH_X1 port map( G => n17734
                           , D => n13184, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_29_3_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_27_3_inst : DLH_X1 port map( G => n17732
                           , D => n13184, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_27_3_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_25_3_inst : DLH_X1 port map( G => n17730
                           , D => n13184, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_25_3_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_23_3_inst : DLH_X1 port map( G => n17728
                           , D => n13184, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_23_3_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_21_3_inst : DLH_X1 port map( G => n17726
                           , D => n13184, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_21_3_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_19_3_inst : DLH_X1 port map( G => n17724
                           , D => n13184, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_19_3_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_17_3_inst : DLH_X1 port map( G => n17722
                           , D => n13184, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_17_3_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_15_3_inst : DLH_X1 port map( G => n17720
                           , D => n13184, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_15_3_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_13_3_inst : DLH_X1 port map( G => n17718
                           , D => n13184, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_13_3_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_11_3_inst : DLH_X1 port map( G => n17716
                           , D => n13184, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_11_3_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_9_3_inst : DLH_X1 port map( G => n17714,
                           D => n13184, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_9_3_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_7_3_inst : DLH_X1 port map( G => n17712,
                           D => n13184, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_7_3_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_5_3_inst : DLH_X1 port map( G => n17710,
                           D => n13184, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_5_3_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_3_3_inst : DLH_X1 port map( G => n17708,
                           D => n13184, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_3_3_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_1_3_inst : DLH_X1 port map( G => n17706,
                           D => n13184, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_1_3_port);
   pipeline_IDEX_Stage_Reg2_out_IDEX_reg_3_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N137, CK => Clk, Q => n13846, QN
                           => n17498);
   pipeline_stageF_PC_reg_PC_out_reg_3_inst : DFFR_X1 port map( D => n3878, CK 
                           => Clk, RN => n17704, Q => n13845, QN => n7658);
   pipeline_IDEX_Stage_Reg1_out_IDEX_reg_3_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N105, CK => Clk, Q => n13844, QN
                           => net214750);
   DataMem_Mem_reg_0_6_inst : DLH_X1 port map( G => n13058, D => DataMem_N1661,
                           Q => DataMem_Mem_0_6_port);
   DataMem_Dataout_reg_6_inst : DLL_X1 port map( D => DataMem_N2179, GN => 
                           n17098, Q => DataMem_N2331);
   pipeline_MEMWB_Stage_Data_to_RF_reg_6_inst : DFF_X1 port map( D => 
                           pipeline_MEMWB_Stage_N17, CK => Clk, Q => 
                           pipeline_data_to_RF_from_WB_6_port, QN => n17318);
   pipeline_RegFile_DEC_WB_RegBank_reg_2_6_inst : DLH_X1 port map( G => n17707,
                           D => n13193, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_2_6_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_4_6_inst : DLH_X1 port map( G => n17709,
                           D => n13193, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_4_6_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_6_6_inst : DLH_X1 port map( G => n17711,
                           D => n13193, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_6_6_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_8_6_inst : DLH_X1 port map( G => n17713,
                           D => n13193, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_8_6_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_10_6_inst : DLH_X1 port map( G => n17715
                           , D => n13193, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_10_6_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_12_6_inst : DLH_X1 port map( G => n17717
                           , D => n13193, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_12_6_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_14_6_inst : DLH_X1 port map( G => n17719
                           , D => n13193, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_14_6_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_16_6_inst : DLH_X1 port map( G => n17721
                           , D => n13193, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_16_6_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_18_6_inst : DLH_X1 port map( G => n17723
                           , D => n13193, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_18_6_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_20_6_inst : DLH_X1 port map( G => n17725
                           , D => n13193, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_20_6_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_22_6_inst : DLH_X1 port map( G => n17727
                           , D => n13193, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_22_6_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_24_6_inst : DLH_X1 port map( G => n17729
                           , D => n13193, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_24_6_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_26_6_inst : DLH_X1 port map( G => n17731
                           , D => n13193, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_26_6_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_28_6_inst : DLH_X1 port map( G => n17733
                           , D => n13193, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_28_6_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_30_6_inst : DLH_X1 port map( G => n17735
                           , D => n13193, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_30_6_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_31_6_inst : DLH_X1 port map( G => n17736
                           , D => n13193, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_31_6_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_29_6_inst : DLH_X1 port map( G => n17734
                           , D => n13193, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_29_6_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_27_6_inst : DLH_X1 port map( G => n17732
                           , D => n13193, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_27_6_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_25_6_inst : DLH_X1 port map( G => n17730
                           , D => n13193, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_25_6_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_23_6_inst : DLH_X1 port map( G => n17728
                           , D => n13193, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_23_6_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_21_6_inst : DLH_X1 port map( G => n17726
                           , D => n13193, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_21_6_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_19_6_inst : DLH_X1 port map( G => n17724
                           , D => n13193, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_19_6_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_17_6_inst : DLH_X1 port map( G => n17722
                           , D => n13193, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_17_6_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_15_6_inst : DLH_X1 port map( G => n17720
                           , D => n13193, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_15_6_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_13_6_inst : DLH_X1 port map( G => n17718
                           , D => n13193, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_13_6_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_11_6_inst : DLH_X1 port map( G => n17716
                           , D => n13193, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_11_6_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_9_6_inst : DLH_X1 port map( G => n17714,
                           D => n13193, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_9_6_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_7_6_inst : DLH_X1 port map( G => n17712,
                           D => n13193, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_7_6_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_5_6_inst : DLH_X1 port map( G => n17710,
                           D => n13193, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_5_6_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_3_6_inst : DLH_X1 port map( G => n17708,
                           D => n13193, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_3_6_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_1_6_inst : DLH_X1 port map( G => n17706,
                           D => n13193, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_1_6_port);
   pipeline_IDEX_Stage_Reg2_out_IDEX_reg_6_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N140, CK => Clk, Q => n13843, QN
                           => n17501);
   pipeline_IDEX_Stage_Reg1_out_IDEX_reg_6_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N108, CK => Clk, Q => n13842, QN
                           => net214749);
   pipeline_EXMEM_stage_ALUres_MEMaddr_out_EXMEM_reg_7_inst : DFF_X1 port map( 
                           D => pipeline_EXMEM_stage_N14, CK => Clk, Q => 
                           pipeline_Alu_Out_Addr_to_mem_7_port, QN => net214748
                           );
   pipeline_MEMWB_Stage_Data_to_RF_reg_7_inst : DFF_X1 port map( D => 
                           pipeline_MEMWB_Stage_N18, CK => Clk, Q => 
                           pipeline_data_to_RF_from_WB_7_port, QN => n17343);
   pipeline_RegFile_DEC_WB_RegBank_reg_2_7_inst : DLH_X1 port map( G => n17707,
                           D => n13196, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_2_7_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_4_7_inst : DLH_X1 port map( G => n17709,
                           D => n13196, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_4_7_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_6_7_inst : DLH_X1 port map( G => n17711,
                           D => n13196, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_6_7_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_8_7_inst : DLH_X1 port map( G => n17713,
                           D => n13196, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_8_7_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_10_7_inst : DLH_X1 port map( G => n17715
                           , D => n13196, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_10_7_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_12_7_inst : DLH_X1 port map( G => n17717
                           , D => n13196, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_12_7_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_14_7_inst : DLH_X1 port map( G => n17719
                           , D => n13196, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_14_7_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_16_7_inst : DLH_X1 port map( G => n17721
                           , D => n13196, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_16_7_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_18_7_inst : DLH_X1 port map( G => n17723
                           , D => n13196, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_18_7_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_20_7_inst : DLH_X1 port map( G => n17725
                           , D => n13196, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_20_7_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_22_7_inst : DLH_X1 port map( G => n17727
                           , D => n13196, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_22_7_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_24_7_inst : DLH_X1 port map( G => n17729
                           , D => n13196, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_24_7_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_26_7_inst : DLH_X1 port map( G => n17731
                           , D => n13196, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_26_7_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_28_7_inst : DLH_X1 port map( G => n17733
                           , D => n13196, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_28_7_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_30_7_inst : DLH_X1 port map( G => n17735
                           , D => n13196, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_30_7_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_31_7_inst : DLH_X1 port map( G => n17736
                           , D => n13196, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_31_7_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_29_7_inst : DLH_X1 port map( G => n17734
                           , D => n13196, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_29_7_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_27_7_inst : DLH_X1 port map( G => n17732
                           , D => n13196, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_27_7_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_25_7_inst : DLH_X1 port map( G => n17730
                           , D => n13196, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_25_7_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_23_7_inst : DLH_X1 port map( G => n17728
                           , D => n13196, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_23_7_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_21_7_inst : DLH_X1 port map( G => n17726
                           , D => n13196, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_21_7_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_19_7_inst : DLH_X1 port map( G => n17724
                           , D => n13196, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_19_7_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_17_7_inst : DLH_X1 port map( G => n17722
                           , D => n13196, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_17_7_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_15_7_inst : DLH_X1 port map( G => n17720
                           , D => n13196, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_15_7_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_13_7_inst : DLH_X1 port map( G => n17718
                           , D => n13196, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_13_7_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_11_7_inst : DLH_X1 port map( G => n17716
                           , D => n13196, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_11_7_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_9_7_inst : DLH_X1 port map( G => n17714,
                           D => n13196, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_9_7_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_7_7_inst : DLH_X1 port map( G => n17712,
                           D => n13196, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_7_7_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_5_7_inst : DLH_X1 port map( G => n17710,
                           D => n13196, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_5_7_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_3_7_inst : DLH_X1 port map( G => n17708,
                           D => n13196, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_3_7_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_1_7_inst : DLH_X1 port map( G => n17706,
                           D => n13196, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_1_7_port);
   pipeline_IDEX_Stage_Reg2_out_IDEX_reg_7_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N141, CK => Clk, Q => n13841, QN
                           => n17502);
   pipeline_stageF_PC_reg_PC_out_reg_7_inst : DFFR_X1 port map( D => n3876, CK 
                           => Clk, RN => n17705, Q => n13840, QN => n7657);
   pipeline_IDEX_Stage_Reg1_out_IDEX_reg_7_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N109, CK => Clk, Q => n13839, QN
                           => net214747);
   DataMem_Mem_reg_7_1_inst : DLH_X1 port map( G => n13079, D => DataMem_N2099,
                           Q => DataMem_Mem_7_1_port);
   DataMem_Mem_reg_6_1_inst : DLH_X1 port map( G => n13076, D => DataMem_N2035,
                           Q => DataMem_Mem_6_1_port);
   DataMem_Mem_reg_5_1_inst : DLH_X1 port map( G => n13073, D => DataMem_N1971,
                           Q => DataMem_Mem_5_1_port);
   DataMem_Mem_reg_4_1_inst : DLH_X1 port map( G => n13070, D => DataMem_N1907,
                           Q => DataMem_Mem_4_1_port);
   DataMem_Mem_reg_3_1_inst : DLH_X1 port map( G => n13067, D => DataMem_N1843,
                           Q => DataMem_Mem_3_1_port);
   DataMem_Mem_reg_2_1_inst : DLH_X1 port map( G => n13064, D => DataMem_N1779,
                           Q => DataMem_Mem_2_1_port);
   DataMem_Mem_reg_1_1_inst : DLH_X1 port map( G => n13061, D => DataMem_N1715,
                           Q => DataMem_Mem_1_1_port);
   pipeline_MEMWB_Stage_Data_to_RF_reg_4_inst : DFF_X1 port map( D => 
                           pipeline_MEMWB_Stage_N15, CK => Clk, Q => 
                           pipeline_data_to_RF_from_WB_4_port, QN => n17320);
   pipeline_RegFile_DEC_WB_RegBank_reg_2_4_inst : DLH_X1 port map( G => n17707,
                           D => n13187, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_2_4_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_4_4_inst : DLH_X1 port map( G => n17709,
                           D => n13187, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_4_4_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_6_4_inst : DLH_X1 port map( G => n17711,
                           D => n13187, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_6_4_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_8_4_inst : DLH_X1 port map( G => n17713,
                           D => n13187, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_8_4_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_10_4_inst : DLH_X1 port map( G => n17715
                           , D => n13187, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_10_4_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_12_4_inst : DLH_X1 port map( G => n17717
                           , D => n13187, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_12_4_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_14_4_inst : DLH_X1 port map( G => n17719
                           , D => n13187, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_14_4_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_16_4_inst : DLH_X1 port map( G => n17721
                           , D => n13187, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_16_4_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_18_4_inst : DLH_X1 port map( G => n17723
                           , D => n13187, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_18_4_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_20_4_inst : DLH_X1 port map( G => n17725
                           , D => n13187, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_20_4_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_22_4_inst : DLH_X1 port map( G => n17727
                           , D => n13187, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_22_4_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_24_4_inst : DLH_X1 port map( G => n17729
                           , D => n13187, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_24_4_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_26_4_inst : DLH_X1 port map( G => n17731
                           , D => n13187, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_26_4_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_28_4_inst : DLH_X1 port map( G => n17733
                           , D => n13187, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_28_4_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_30_4_inst : DLH_X1 port map( G => n17735
                           , D => n13187, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_30_4_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_31_4_inst : DLH_X1 port map( G => n17736
                           , D => n13187, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_31_4_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_29_4_inst : DLH_X1 port map( G => n17734
                           , D => n13187, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_29_4_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_27_4_inst : DLH_X1 port map( G => n17732
                           , D => n13187, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_27_4_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_25_4_inst : DLH_X1 port map( G => n17730
                           , D => n13187, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_25_4_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_23_4_inst : DLH_X1 port map( G => n17728
                           , D => n13187, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_23_4_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_21_4_inst : DLH_X1 port map( G => n17726
                           , D => n13187, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_21_4_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_19_4_inst : DLH_X1 port map( G => n17724
                           , D => n13187, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_19_4_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_17_4_inst : DLH_X1 port map( G => n17722
                           , D => n13187, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_17_4_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_15_4_inst : DLH_X1 port map( G => n17720
                           , D => n13187, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_15_4_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_13_4_inst : DLH_X1 port map( G => n17718
                           , D => n13187, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_13_4_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_11_4_inst : DLH_X1 port map( G => n17716
                           , D => n13187, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_11_4_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_9_4_inst : DLH_X1 port map( G => n17714,
                           D => n13187, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_9_4_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_7_4_inst : DLH_X1 port map( G => n17712,
                           D => n13187, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_7_4_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_5_4_inst : DLH_X1 port map( G => n17710,
                           D => n13187, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_5_4_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_3_4_inst : DLH_X1 port map( G => n17708,
                           D => n13187, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_3_4_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_1_4_inst : DLH_X1 port map( G => n17706,
                           D => n13187, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_1_4_port);
   pipeline_IDEX_Stage_Reg2_out_IDEX_reg_4_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N138, CK => Clk, Q => n13838, QN
                           => n17499);
   pipeline_stageF_PC_reg_PC_out_reg_4_inst : DFFR_X1 port map( D => n3874, CK 
                           => Clk, RN => n17704, Q => n13837, QN => n7656);
   pipeline_IDEX_Stage_Reg1_out_IDEX_reg_4_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N106, CK => Clk, Q => n13836, QN
                           => net214746);
   pipeline_EXMEM_stage_DataToMem_out_EXMEM_reg_4_inst : DFF_X1 port map( D => 
                           pipeline_EXMEM_stage_N43, CK => Clk, Q => n13835, QN
                           => net214745);
   DataMem_Mem_reg_7_4_inst : DLH_X1 port map( G => n13079, D => DataMem_N2105,
                           Q => DataMem_Mem_7_4_port);
   DataMem_Mem_reg_6_4_inst : DLH_X1 port map( G => n13076, D => DataMem_N2041,
                           Q => DataMem_Mem_6_4_port);
   DataMem_Mem_reg_5_4_inst : DLH_X1 port map( G => n13073, D => DataMem_N1977,
                           Q => DataMem_Mem_5_4_port);
   DataMem_Mem_reg_4_4_inst : DLH_X1 port map( G => n13070, D => DataMem_N1913,
                           Q => DataMem_Mem_4_4_port);
   DataMem_Mem_reg_3_4_inst : DLH_X1 port map( G => n13067, D => DataMem_N1849,
                           Q => DataMem_Mem_3_4_port);
   DataMem_Mem_reg_2_4_inst : DLH_X1 port map( G => n13064, D => DataMem_N1785,
                           Q => DataMem_Mem_2_4_port);
   DataMem_Mem_reg_1_4_inst : DLH_X1 port map( G => n13061, D => DataMem_N1721,
                           Q => DataMem_Mem_1_4_port);
   DataMem_Mem_reg_0_4_inst : DLH_X1 port map( G => n13058, D => DataMem_N1657,
                           Q => DataMem_Mem_0_4_port);
   DataMem_Dataout_reg_4_inst : DLL_X1 port map( D => DataMem_N2173, GN => 
                           n17098, Q => DataMem_N2337);
   pipeline_MEMWB_Stage_Data_to_RF_reg_5_inst : DFF_X1 port map( D => 
                           pipeline_MEMWB_Stage_N16, CK => Clk, Q => 
                           pipeline_data_to_RF_from_WB_5_port, QN => n17308);
   pipeline_RegFile_DEC_WB_RegBank_reg_2_5_inst : DLH_X1 port map( G => n13169,
                           D => n13190, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_2_5_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_4_5_inst : DLH_X1 port map( G => n13163,
                           D => n13190, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_4_5_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_6_5_inst : DLH_X1 port map( G => n13157,
                           D => n13190, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_6_5_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_8_5_inst : DLH_X1 port map( G => n13151,
                           D => n13190, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_8_5_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_10_5_inst : DLH_X1 port map( G => n13145
                           , D => n13190, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_10_5_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_12_5_inst : DLH_X1 port map( G => n13139
                           , D => n13190, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_12_5_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_14_5_inst : DLH_X1 port map( G => n13133
                           , D => n13190, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_14_5_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_16_5_inst : DLH_X1 port map( G => n13127
                           , D => n13190, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_16_5_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_18_5_inst : DLH_X1 port map( G => n13121
                           , D => n13190, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_18_5_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_20_5_inst : DLH_X1 port map( G => n13115
                           , D => n13190, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_20_5_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_22_5_inst : DLH_X1 port map( G => n13109
                           , D => n13190, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_22_5_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_24_5_inst : DLH_X1 port map( G => n13103
                           , D => n13190, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_24_5_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_26_5_inst : DLH_X1 port map( G => n13097
                           , D => n13190, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_26_5_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_28_5_inst : DLH_X1 port map( G => n13091
                           , D => n13190, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_28_5_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_30_5_inst : DLH_X1 port map( G => n13085
                           , D => n13190, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_30_5_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_31_5_inst : DLH_X1 port map( G => n13082
                           , D => n13190, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_31_5_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_29_5_inst : DLH_X1 port map( G => n13088
                           , D => n13190, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_29_5_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_27_5_inst : DLH_X1 port map( G => n13094
                           , D => n13190, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_27_5_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_25_5_inst : DLH_X1 port map( G => n13100
                           , D => n13190, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_25_5_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_23_5_inst : DLH_X1 port map( G => n13106
                           , D => n13190, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_23_5_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_21_5_inst : DLH_X1 port map( G => n13112
                           , D => n13190, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_21_5_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_19_5_inst : DLH_X1 port map( G => n13118
                           , D => n13190, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_19_5_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_17_5_inst : DLH_X1 port map( G => n13124
                           , D => n13190, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_17_5_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_15_5_inst : DLH_X1 port map( G => n13130
                           , D => n13190, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_15_5_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_13_5_inst : DLH_X1 port map( G => n13136
                           , D => n13190, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_13_5_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_11_5_inst : DLH_X1 port map( G => n13142
                           , D => n13190, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_11_5_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_9_5_inst : DLH_X1 port map( G => n13148,
                           D => n13190, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_9_5_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_7_5_inst : DLH_X1 port map( G => n13154,
                           D => n13190, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_7_5_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_5_5_inst : DLH_X1 port map( G => n13160,
                           D => n13190, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_5_5_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_3_5_inst : DLH_X1 port map( G => n13166,
                           D => n13190, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_3_5_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_1_5_inst : DLH_X1 port map( G => n13172,
                           D => n13190, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_1_5_port);
   pipeline_IDEX_Stage_Reg2_out_IDEX_reg_5_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N139, CK => Clk, Q => n13834, QN
                           => n17500);
   pipeline_stageF_PC_reg_PC_out_reg_5_inst : DFFR_X1 port map( D => n3872, CK 
                           => Clk, RN => n17705, Q => n13833, QN => n7655);
   pipeline_IDEX_Stage_Reg1_out_IDEX_reg_5_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N107, CK => Clk, Q => n13832, QN
                           => net214744);
   pipeline_EXMEM_stage_DataToMem_out_EXMEM_reg_5_inst : DFF_X1 port map( D => 
                           pipeline_EXMEM_stage_N44, CK => Clk, Q => n13831, QN
                           => net214743);
   DataMem_Mem_reg_7_5_inst : DLH_X1 port map( G => n13079, D => DataMem_N2107,
                           Q => DataMem_Mem_7_5_port);
   DataMem_Mem_reg_6_5_inst : DLH_X1 port map( G => n13076, D => DataMem_N2043,
                           Q => DataMem_Mem_6_5_port);
   DataMem_Mem_reg_5_5_inst : DLH_X1 port map( G => n13073, D => DataMem_N1979,
                           Q => DataMem_Mem_5_5_port);
   DataMem_Mem_reg_4_5_inst : DLH_X1 port map( G => n13070, D => DataMem_N1915,
                           Q => DataMem_Mem_4_5_port);
   DataMem_Mem_reg_3_5_inst : DLH_X1 port map( G => n13067, D => DataMem_N1851,
                           Q => DataMem_Mem_3_5_port);
   DataMem_Mem_reg_2_5_inst : DLH_X1 port map( G => n13064, D => DataMem_N1787,
                           Q => DataMem_Mem_2_5_port);
   DataMem_Mem_reg_1_5_inst : DLH_X1 port map( G => n13061, D => DataMem_N1723,
                           Q => DataMem_Mem_1_5_port);
   DataMem_Mem_reg_0_5_inst : DLH_X1 port map( G => n13058, D => DataMem_N1659,
                           Q => DataMem_Mem_0_5_port);
   DataMem_Dataout_reg_5_inst : DLL_X1 port map( D => DataMem_N2176, GN => 
                           n17098, Q => DataMem_N2334);
   pipeline_EXMEM_stage_DataToMem_out_EXMEM_reg_7_inst : DFF_X1 port map( D => 
                           pipeline_EXMEM_stage_N46, CK => Clk, Q => n13830, QN
                           => net214742);
   DataMem_Mem_reg_7_7_inst : DLH_X1 port map( G => n13079, D => DataMem_N2111,
                           Q => DataMem_Mem_7_7_port);
   DataMem_Mem_reg_6_7_inst : DLH_X1 port map( G => n13076, D => DataMem_N2047,
                           Q => DataMem_Mem_6_7_port);
   DataMem_Mem_reg_5_7_inst : DLH_X1 port map( G => n13073, D => DataMem_N1983,
                           Q => DataMem_Mem_5_7_port);
   DataMem_Mem_reg_4_7_inst : DLH_X1 port map( G => n13070, D => DataMem_N1919,
                           Q => DataMem_Mem_4_7_port);
   DataMem_Mem_reg_3_7_inst : DLH_X1 port map( G => n13067, D => DataMem_N1855,
                           Q => DataMem_Mem_3_7_port);
   DataMem_Mem_reg_2_7_inst : DLH_X1 port map( G => n13064, D => DataMem_N1791,
                           Q => DataMem_Mem_2_7_port);
   DataMem_Mem_reg_1_7_inst : DLH_X1 port map( G => n13061, D => DataMem_N1727,
                           Q => DataMem_Mem_1_7_port);
   DataMem_Mem_reg_0_7_inst : DLH_X1 port map( G => n13058, D => DataMem_N1663,
                           Q => DataMem_Mem_0_7_port);
   DataMem_Dataout_reg_7_inst : DLL_X1 port map( D => DataMem_N2182, GN => 
                           n17098, Q => DataMem_N2328);
   pipeline_stageF_PC_reg_PC_out_reg_6_inst : DFFR_X1 port map( D => n3870, CK 
                           => Clk, RN => n17705, Q => n13829, QN => n7654);
   pipeline_EXMEM_stage_DataToMem_out_EXMEM_reg_6_inst : DFF_X1 port map( D => 
                           pipeline_EXMEM_stage_N45, CK => Clk, Q => n13828, QN
                           => net214741);
   DataMem_Mem_reg_7_6_inst : DLH_X1 port map( G => n13079, D => DataMem_N2109,
                           Q => DataMem_Mem_7_6_port);
   DataMem_Mem_reg_6_6_inst : DLH_X1 port map( G => n13076, D => DataMem_N2045,
                           Q => DataMem_Mem_6_6_port);
   DataMem_Mem_reg_5_6_inst : DLH_X1 port map( G => n13073, D => DataMem_N1981,
                           Q => DataMem_Mem_5_6_port);
   DataMem_Mem_reg_4_6_inst : DLH_X1 port map( G => n13070, D => DataMem_N1917,
                           Q => DataMem_Mem_4_6_port);
   DataMem_Mem_reg_3_6_inst : DLH_X1 port map( G => n13067, D => DataMem_N1853,
                           Q => DataMem_Mem_3_6_port);
   DataMem_Mem_reg_2_6_inst : DLH_X1 port map( G => n13064, D => DataMem_N1789,
                           Q => DataMem_Mem_2_6_port);
   DataMem_Mem_reg_1_6_inst : DLH_X1 port map( G => n13061, D => DataMem_N1725,
                           Q => DataMem_Mem_1_6_port);
   DataMem_Mem_reg_0_10_inst : DLH_X1 port map( G => n13058, D => DataMem_N1669
                           , Q => DataMem_Mem_0_10_port);
   DataMem_Dataout_reg_10_inst : DLL_X1 port map( D => DataMem_N2191, GN => 
                           n13055, Q => DataMem_N2319);
   pipeline_MEMWB_Stage_Data_to_RF_reg_10_inst : DFF_X1 port map( D => 
                           pipeline_MEMWB_Stage_N21, CK => Clk, Q => 
                           pipeline_data_to_RF_from_WB_10_port, QN => n17307);
   pipeline_RegFile_DEC_WB_RegBank_reg_2_10_inst : DLH_X1 port map( G => n13169
                           , D => n13205, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_2_10_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_4_10_inst : DLH_X1 port map( G => n13163
                           , D => n13205, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_4_10_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_6_10_inst : DLH_X1 port map( G => n13157
                           , D => n13205, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_6_10_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_8_10_inst : DLH_X1 port map( G => n13151
                           , D => n13205, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_8_10_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_10_10_inst : DLH_X1 port map( G => 
                           n13145, D => n13205, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_10_10_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_12_10_inst : DLH_X1 port map( G => 
                           n13139, D => n13205, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_12_10_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_14_10_inst : DLH_X1 port map( G => 
                           n13133, D => n13205, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_14_10_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_16_10_inst : DLH_X1 port map( G => 
                           n13127, D => n13205, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_16_10_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_18_10_inst : DLH_X1 port map( G => 
                           n13121, D => n13205, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_18_10_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_20_10_inst : DLH_X1 port map( G => 
                           n13115, D => n13205, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_20_10_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_22_10_inst : DLH_X1 port map( G => 
                           n13109, D => n13205, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_22_10_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_24_10_inst : DLH_X1 port map( G => 
                           n13103, D => n13205, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_24_10_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_26_10_inst : DLH_X1 port map( G => 
                           n13097, D => n13205, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_26_10_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_28_10_inst : DLH_X1 port map( G => 
                           n13091, D => n13205, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_28_10_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_30_10_inst : DLH_X1 port map( G => 
                           n13085, D => n13205, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_30_10_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_31_10_inst : DLH_X1 port map( G => 
                           n13082, D => n13205, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_31_10_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_29_10_inst : DLH_X1 port map( G => 
                           n13088, D => n13205, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_29_10_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_27_10_inst : DLH_X1 port map( G => 
                           n13094, D => n13205, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_27_10_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_25_10_inst : DLH_X1 port map( G => 
                           n13100, D => n13205, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_25_10_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_23_10_inst : DLH_X1 port map( G => 
                           n13106, D => n13205, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_23_10_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_21_10_inst : DLH_X1 port map( G => 
                           n13112, D => n13205, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_21_10_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_19_10_inst : DLH_X1 port map( G => 
                           n13118, D => n13205, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_19_10_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_17_10_inst : DLH_X1 port map( G => 
                           n13124, D => n13205, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_17_10_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_15_10_inst : DLH_X1 port map( G => 
                           n13130, D => n13205, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_15_10_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_13_10_inst : DLH_X1 port map( G => 
                           n13136, D => n13205, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_13_10_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_11_10_inst : DLH_X1 port map( G => 
                           n13142, D => n13205, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_11_10_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_9_10_inst : DLH_X1 port map( G => n13148
                           , D => n13205, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_9_10_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_7_10_inst : DLH_X1 port map( G => n13154
                           , D => n13205, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_7_10_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_5_10_inst : DLH_X1 port map( G => n13160
                           , D => n13205, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_5_10_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_3_10_inst : DLH_X1 port map( G => n13166
                           , D => n13205, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_3_10_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_1_10_inst : DLH_X1 port map( G => n13172
                           , D => n13205, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_1_10_port);
   pipeline_IDEX_Stage_Reg2_out_IDEX_reg_10_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N144, CK => Clk, Q => n13827, QN
                           => n17505);
   pipeline_IDEX_Stage_Reg1_out_IDEX_reg_10_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N112, CK => Clk, Q => n13826, QN
                           => net214740);
   pipeline_MEMWB_Stage_Data_to_RF_reg_11_inst : DFF_X1 port map( D => 
                           pipeline_MEMWB_Stage_N22, CK => Clk, Q => 
                           pipeline_data_to_RF_from_WB_11_port, QN => n17319);
   pipeline_RegFile_DEC_WB_RegBank_reg_2_11_inst : DLH_X1 port map( G => n17707
                           , D => n13208, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_2_11_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_4_11_inst : DLH_X1 port map( G => n17709
                           , D => n13208, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_4_11_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_6_11_inst : DLH_X1 port map( G => n17711
                           , D => n13208, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_6_11_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_8_11_inst : DLH_X1 port map( G => n17713
                           , D => n13208, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_8_11_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_10_11_inst : DLH_X1 port map( G => 
                           n17715, D => n13208, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_10_11_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_12_11_inst : DLH_X1 port map( G => 
                           n17717, D => n13208, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_12_11_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_14_11_inst : DLH_X1 port map( G => 
                           n17719, D => n13208, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_14_11_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_16_11_inst : DLH_X1 port map( G => 
                           n17721, D => n13208, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_16_11_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_18_11_inst : DLH_X1 port map( G => 
                           n17723, D => n13208, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_18_11_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_20_11_inst : DLH_X1 port map( G => 
                           n17725, D => n13208, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_20_11_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_22_11_inst : DLH_X1 port map( G => 
                           n17727, D => n13208, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_22_11_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_24_11_inst : DLH_X1 port map( G => 
                           n17729, D => n13208, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_24_11_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_26_11_inst : DLH_X1 port map( G => 
                           n17731, D => n13208, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_26_11_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_28_11_inst : DLH_X1 port map( G => 
                           n17733, D => n13208, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_28_11_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_30_11_inst : DLH_X1 port map( G => 
                           n17735, D => n13208, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_30_11_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_31_11_inst : DLH_X1 port map( G => 
                           n17736, D => n13208, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_31_11_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_29_11_inst : DLH_X1 port map( G => 
                           n17734, D => n13208, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_29_11_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_27_11_inst : DLH_X1 port map( G => 
                           n17732, D => n13208, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_27_11_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_25_11_inst : DLH_X1 port map( G => 
                           n17730, D => n13208, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_25_11_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_23_11_inst : DLH_X1 port map( G => 
                           n17728, D => n13208, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_23_11_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_21_11_inst : DLH_X1 port map( G => 
                           n17726, D => n13208, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_21_11_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_19_11_inst : DLH_X1 port map( G => 
                           n17724, D => n13208, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_19_11_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_17_11_inst : DLH_X1 port map( G => 
                           n17722, D => n13208, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_17_11_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_15_11_inst : DLH_X1 port map( G => 
                           n17720, D => n13208, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_15_11_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_13_11_inst : DLH_X1 port map( G => 
                           n17718, D => n13208, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_13_11_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_11_11_inst : DLH_X1 port map( G => 
                           n17716, D => n13208, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_11_11_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_9_11_inst : DLH_X1 port map( G => n17714
                           , D => n13208, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_9_11_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_7_11_inst : DLH_X1 port map( G => n17712
                           , D => n13208, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_7_11_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_5_11_inst : DLH_X1 port map( G => n17710
                           , D => n13208, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_5_11_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_3_11_inst : DLH_X1 port map( G => n17708
                           , D => n13208, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_3_11_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_1_11_inst : DLH_X1 port map( G => n17706
                           , D => n13208, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_1_11_port);
   pipeline_IDEX_Stage_Reg2_out_IDEX_reg_11_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N145, CK => Clk, Q => n13825, QN
                           => n17506);
   pipeline_stageF_PC_reg_PC_out_reg_11_inst : DFFR_X1 port map( D => n3868, CK
                           => Clk, RN => n17704, Q => n13824, QN => n7653);
   pipeline_IDEX_Stage_Reg1_out_IDEX_reg_11_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N113, CK => Clk, Q => n13823, QN
                           => net214739);
   pipeline_MEMWB_Stage_Data_to_RF_reg_9_inst : DFF_X1 port map( D => 
                           pipeline_MEMWB_Stage_N20, CK => Clk, Q => 
                           pipeline_data_to_RF_from_WB_9_port, QN => n17305);
   pipeline_RegFile_DEC_WB_RegBank_reg_2_9_inst : DLH_X1 port map( G => n13169,
                           D => n13202, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_2_9_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_4_9_inst : DLH_X1 port map( G => n13163,
                           D => n13202, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_4_9_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_6_9_inst : DLH_X1 port map( G => n13157,
                           D => n13202, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_6_9_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_8_9_inst : DLH_X1 port map( G => n13151,
                           D => n13202, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_8_9_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_10_9_inst : DLH_X1 port map( G => n13145
                           , D => n13202, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_10_9_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_12_9_inst : DLH_X1 port map( G => n13139
                           , D => n13202, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_12_9_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_14_9_inst : DLH_X1 port map( G => n13133
                           , D => n13202, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_14_9_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_16_9_inst : DLH_X1 port map( G => n13127
                           , D => n13202, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_16_9_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_18_9_inst : DLH_X1 port map( G => n13121
                           , D => n13202, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_18_9_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_20_9_inst : DLH_X1 port map( G => n13115
                           , D => n13202, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_20_9_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_22_9_inst : DLH_X1 port map( G => n13109
                           , D => n13202, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_22_9_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_24_9_inst : DLH_X1 port map( G => n13103
                           , D => n13202, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_24_9_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_26_9_inst : DLH_X1 port map( G => n13097
                           , D => n13202, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_26_9_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_28_9_inst : DLH_X1 port map( G => n13091
                           , D => n13202, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_28_9_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_30_9_inst : DLH_X1 port map( G => n13085
                           , D => n13202, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_30_9_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_31_9_inst : DLH_X1 port map( G => n13082
                           , D => n13202, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_31_9_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_29_9_inst : DLH_X1 port map( G => n13088
                           , D => n13202, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_29_9_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_27_9_inst : DLH_X1 port map( G => n13094
                           , D => n13202, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_27_9_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_25_9_inst : DLH_X1 port map( G => n13100
                           , D => n13202, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_25_9_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_23_9_inst : DLH_X1 port map( G => n13106
                           , D => n13202, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_23_9_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_21_9_inst : DLH_X1 port map( G => n13112
                           , D => n13202, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_21_9_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_19_9_inst : DLH_X1 port map( G => n13118
                           , D => n13202, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_19_9_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_17_9_inst : DLH_X1 port map( G => n13124
                           , D => n13202, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_17_9_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_15_9_inst : DLH_X1 port map( G => n13130
                           , D => n13202, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_15_9_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_13_9_inst : DLH_X1 port map( G => n13136
                           , D => n13202, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_13_9_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_11_9_inst : DLH_X1 port map( G => n13142
                           , D => n13202, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_11_9_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_9_9_inst : DLH_X1 port map( G => n13148,
                           D => n13202, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_9_9_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_7_9_inst : DLH_X1 port map( G => n13154,
                           D => n13202, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_7_9_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_5_9_inst : DLH_X1 port map( G => n13160,
                           D => n13202, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_5_9_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_3_9_inst : DLH_X1 port map( G => n13166,
                           D => n13202, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_3_9_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_1_9_inst : DLH_X1 port map( G => n13172,
                           D => n13202, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_1_9_port);
   pipeline_IDEX_Stage_Reg2_out_IDEX_reg_9_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N143, CK => Clk, Q => n13822, QN
                           => n17504);
   pipeline_stageF_PC_reg_PC_out_reg_9_inst : DFFR_X1 port map( D => n3866, CK 
                           => Clk, RN => n17704, Q => n13821, QN => n7652);
   pipeline_IDEX_Stage_Reg1_out_IDEX_reg_9_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N111, CK => Clk, Q => n13820, QN
                           => net214738);
   pipeline_EXMEM_stage_DataToMem_out_EXMEM_reg_9_inst : DFF_X1 port map( D => 
                           pipeline_EXMEM_stage_N48, CK => Clk, Q => n13819, QN
                           => net214737);
   DataMem_Mem_reg_7_9_inst : DLH_X1 port map( G => n13079, D => DataMem_N2115,
                           Q => DataMem_Mem_7_9_port);
   DataMem_Mem_reg_6_9_inst : DLH_X1 port map( G => n13076, D => DataMem_N2051,
                           Q => DataMem_Mem_6_9_port);
   DataMem_Mem_reg_5_9_inst : DLH_X1 port map( G => n13073, D => DataMem_N1987,
                           Q => DataMem_Mem_5_9_port);
   DataMem_Mem_reg_4_9_inst : DLH_X1 port map( G => n13070, D => DataMem_N1923,
                           Q => DataMem_Mem_4_9_port);
   DataMem_Mem_reg_3_9_inst : DLH_X1 port map( G => n13067, D => DataMem_N1859,
                           Q => DataMem_Mem_3_9_port);
   DataMem_Mem_reg_2_9_inst : DLH_X1 port map( G => n13064, D => DataMem_N1795,
                           Q => DataMem_Mem_2_9_port);
   DataMem_Mem_reg_1_9_inst : DLH_X1 port map( G => n13061, D => DataMem_N1731,
                           Q => DataMem_Mem_1_9_port);
   DataMem_Mem_reg_0_9_inst : DLH_X1 port map( G => n13058, D => DataMem_N1667,
                           Q => DataMem_Mem_0_9_port);
   DataMem_Dataout_reg_9_inst : DLL_X1 port map( D => DataMem_N2188, GN => 
                           n13055, Q => DataMem_N2322);
   pipeline_EXMEM_stage_DataToMem_out_EXMEM_reg_11_inst : DFF_X1 port map( D =>
                           pipeline_EXMEM_stage_N50, CK => Clk, Q => n13818, QN
                           => net214736);
   DataMem_Mem_reg_7_11_inst : DLH_X1 port map( G => n13079, D => DataMem_N2119
                           , Q => DataMem_Mem_7_11_port);
   DataMem_Mem_reg_6_11_inst : DLH_X1 port map( G => n13076, D => DataMem_N2055
                           , Q => DataMem_Mem_6_11_port);
   DataMem_Mem_reg_5_11_inst : DLH_X1 port map( G => n13073, D => DataMem_N1991
                           , Q => DataMem_Mem_5_11_port);
   DataMem_Mem_reg_4_11_inst : DLH_X1 port map( G => n13070, D => DataMem_N1927
                           , Q => DataMem_Mem_4_11_port);
   DataMem_Mem_reg_3_11_inst : DLH_X1 port map( G => n13067, D => DataMem_N1863
                           , Q => DataMem_Mem_3_11_port);
   DataMem_Mem_reg_2_11_inst : DLH_X1 port map( G => n13064, D => DataMem_N1799
                           , Q => DataMem_Mem_2_11_port);
   DataMem_Mem_reg_1_11_inst : DLH_X1 port map( G => n13061, D => DataMem_N1735
                           , Q => DataMem_Mem_1_11_port);
   DataMem_Mem_reg_0_11_inst : DLH_X1 port map( G => n13058, D => DataMem_N1671
                           , Q => DataMem_Mem_0_11_port);
   DataMem_Dataout_reg_11_inst : DLL_X1 port map( D => DataMem_N2194, GN => 
                           n13055, Q => DataMem_N2316);
   pipeline_stageF_PC_reg_PC_out_reg_10_inst : DFFR_X1 port map( D => n3864, CK
                           => Clk, RN => n17705, Q => n13817, QN => n7651);
   pipeline_EXMEM_stage_DataToMem_out_EXMEM_reg_10_inst : DFF_X1 port map( D =>
                           pipeline_EXMEM_stage_N49, CK => Clk, Q => n13816, QN
                           => net214735);
   DataMem_Mem_reg_7_10_inst : DLH_X1 port map( G => n13079, D => DataMem_N2117
                           , Q => DataMem_Mem_7_10_port);
   DataMem_Mem_reg_6_10_inst : DLH_X1 port map( G => n13076, D => DataMem_N2053
                           , Q => DataMem_Mem_6_10_port);
   DataMem_Mem_reg_5_10_inst : DLH_X1 port map( G => n13073, D => DataMem_N1989
                           , Q => DataMem_Mem_5_10_port);
   DataMem_Mem_reg_4_10_inst : DLH_X1 port map( G => n13070, D => DataMem_N1925
                           , Q => DataMem_Mem_4_10_port);
   DataMem_Mem_reg_3_10_inst : DLH_X1 port map( G => n13067, D => DataMem_N1861
                           , Q => DataMem_Mem_3_10_port);
   DataMem_Mem_reg_2_10_inst : DLH_X1 port map( G => n13064, D => DataMem_N1797
                           , Q => DataMem_Mem_2_10_port);
   DataMem_Mem_reg_1_10_inst : DLH_X1 port map( G => n13061, D => DataMem_N1733
                           , Q => DataMem_Mem_1_10_port);
   DataMem_Mem_reg_0_12_inst : DLH_X1 port map( G => n13058, D => DataMem_N1673
                           , Q => DataMem_Mem_0_12_port);
   DataMem_Dataout_reg_12_inst : DLL_X1 port map( D => DataMem_N2197, GN => 
                           n13055, Q => DataMem_N2313);
   pipeline_MEMWB_Stage_Data_to_RF_reg_12_inst : DFF_X1 port map( D => 
                           pipeline_MEMWB_Stage_N23, CK => Clk, Q => 
                           pipeline_data_to_RF_from_WB_12_port, QN => n17395);
   pipeline_RegFile_DEC_WB_RegBank_reg_2_12_inst : DLH_X1 port map( G => n13169
                           , D => n13211, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_2_12_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_4_12_inst : DLH_X1 port map( G => n13163
                           , D => n13211, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_4_12_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_6_12_inst : DLH_X1 port map( G => n13157
                           , D => n13211, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_6_12_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_8_12_inst : DLH_X1 port map( G => n13151
                           , D => n13211, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_8_12_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_10_12_inst : DLH_X1 port map( G => 
                           n13145, D => n13211, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_10_12_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_12_12_inst : DLH_X1 port map( G => 
                           n13139, D => n13211, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_12_12_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_14_12_inst : DLH_X1 port map( G => 
                           n13133, D => n13211, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_14_12_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_16_12_inst : DLH_X1 port map( G => 
                           n13127, D => n13211, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_16_12_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_18_12_inst : DLH_X1 port map( G => 
                           n13121, D => n13211, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_18_12_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_20_12_inst : DLH_X1 port map( G => 
                           n13115, D => n13211, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_20_12_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_22_12_inst : DLH_X1 port map( G => 
                           n13109, D => n13211, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_22_12_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_24_12_inst : DLH_X1 port map( G => 
                           n13103, D => n13211, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_24_12_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_26_12_inst : DLH_X1 port map( G => 
                           n13097, D => n13211, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_26_12_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_28_12_inst : DLH_X1 port map( G => 
                           n13091, D => n13211, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_28_12_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_30_12_inst : DLH_X1 port map( G => 
                           n13085, D => n13211, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_30_12_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_31_12_inst : DLH_X1 port map( G => 
                           n13082, D => n13211, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_31_12_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_29_12_inst : DLH_X1 port map( G => 
                           n13088, D => n13211, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_29_12_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_27_12_inst : DLH_X1 port map( G => 
                           n13094, D => n13211, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_27_12_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_25_12_inst : DLH_X1 port map( G => 
                           n13100, D => n13211, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_25_12_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_23_12_inst : DLH_X1 port map( G => 
                           n13106, D => n13211, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_23_12_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_21_12_inst : DLH_X1 port map( G => 
                           n13112, D => n13211, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_21_12_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_19_12_inst : DLH_X1 port map( G => 
                           n13118, D => n13211, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_19_12_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_17_12_inst : DLH_X1 port map( G => 
                           n13124, D => n13211, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_17_12_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_15_12_inst : DLH_X1 port map( G => 
                           n13130, D => n13211, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_15_12_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_13_12_inst : DLH_X1 port map( G => 
                           n13136, D => n13211, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_13_12_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_11_12_inst : DLH_X1 port map( G => 
                           n13142, D => n13211, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_11_12_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_9_12_inst : DLH_X1 port map( G => n13148
                           , D => n13211, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_9_12_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_7_12_inst : DLH_X1 port map( G => n13154
                           , D => n13211, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_7_12_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_5_12_inst : DLH_X1 port map( G => n13160
                           , D => n13211, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_5_12_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_3_12_inst : DLH_X1 port map( G => n13166
                           , D => n13211, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_3_12_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_1_12_inst : DLH_X1 port map( G => n13172
                           , D => n13211, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_1_12_port);
   pipeline_IDEX_Stage_Reg2_out_IDEX_reg_12_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N146, CK => Clk, Q => n13815, QN
                           => n17507);
   pipeline_IDEX_Stage_Reg1_out_IDEX_reg_12_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N114, CK => Clk, Q => n13814, QN
                           => net214734);
   pipeline_EXMEM_stage_ALUres_MEMaddr_out_EXMEM_reg_12_inst : DFF_X1 port map(
                           D => pipeline_EXMEM_stage_N19, CK => Clk, Q => 
                           pipeline_Alu_Out_Addr_to_mem_12_port, QN => 
                           net214733);
   pipeline_stageF_PC_reg_PC_out_reg_12_inst : DFFR_X1 port map( D => n3862, CK
                           => Clk, RN => n17705, Q => n13813, QN => n7650);
   pipeline_EXMEM_stage_DataToMem_out_EXMEM_reg_12_inst : DFF_X1 port map( D =>
                           pipeline_EXMEM_stage_N51, CK => Clk, Q => n13812, QN
                           => net214732);
   DataMem_Mem_reg_7_12_inst : DLH_X1 port map( G => n13079, D => DataMem_N2121
                           , Q => DataMem_Mem_7_12_port);
   DataMem_Mem_reg_6_12_inst : DLH_X1 port map( G => n13076, D => DataMem_N2057
                           , Q => DataMem_Mem_6_12_port);
   DataMem_Mem_reg_5_12_inst : DLH_X1 port map( G => n13073, D => DataMem_N1993
                           , Q => DataMem_Mem_5_12_port);
   DataMem_Mem_reg_4_12_inst : DLH_X1 port map( G => n13070, D => DataMem_N1929
                           , Q => DataMem_Mem_4_12_port);
   DataMem_Mem_reg_3_12_inst : DLH_X1 port map( G => n13067, D => DataMem_N1865
                           , Q => DataMem_Mem_3_12_port);
   DataMem_Mem_reg_2_12_inst : DLH_X1 port map( G => n13064, D => DataMem_N1801
                           , Q => DataMem_Mem_2_12_port);
   DataMem_Mem_reg_1_12_inst : DLH_X1 port map( G => n13061, D => DataMem_N1737
                           , Q => DataMem_Mem_1_12_port);
   pipeline_MEMWB_Stage_Data_to_RF_reg_2_inst : DFF_X1 port map( D => 
                           pipeline_MEMWB_Stage_N13, CK => Clk, Q => 
                           pipeline_data_to_RF_from_WB_2_port, QN => n17369);
   pipeline_RegFile_DEC_WB_RegBank_reg_2_2_inst : DLH_X1 port map( G => n17707,
                           D => n13181, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_2_2_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_4_2_inst : DLH_X1 port map( G => n17709,
                           D => n13181, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_4_2_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_6_2_inst : DLH_X1 port map( G => n17711,
                           D => n13181, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_6_2_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_8_2_inst : DLH_X1 port map( G => n17713,
                           D => n13181, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_8_2_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_10_2_inst : DLH_X1 port map( G => n17715
                           , D => n13181, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_10_2_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_12_2_inst : DLH_X1 port map( G => n17717
                           , D => n13181, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_12_2_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_14_2_inst : DLH_X1 port map( G => n17719
                           , D => n13181, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_14_2_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_16_2_inst : DLH_X1 port map( G => n17721
                           , D => n13181, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_16_2_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_18_2_inst : DLH_X1 port map( G => n17723
                           , D => n13181, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_18_2_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_20_2_inst : DLH_X1 port map( G => n17725
                           , D => n13181, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_20_2_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_22_2_inst : DLH_X1 port map( G => n17727
                           , D => n13181, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_22_2_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_24_2_inst : DLH_X1 port map( G => n17729
                           , D => n13181, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_24_2_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_26_2_inst : DLH_X1 port map( G => n17731
                           , D => n13181, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_26_2_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_28_2_inst : DLH_X1 port map( G => n17733
                           , D => n13181, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_28_2_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_30_2_inst : DLH_X1 port map( G => n17735
                           , D => n13181, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_30_2_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_31_2_inst : DLH_X1 port map( G => n17736
                           , D => n13181, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_31_2_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_29_2_inst : DLH_X1 port map( G => n17734
                           , D => n13181, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_29_2_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_27_2_inst : DLH_X1 port map( G => n17732
                           , D => n13181, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_27_2_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_25_2_inst : DLH_X1 port map( G => n17730
                           , D => n13181, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_25_2_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_23_2_inst : DLH_X1 port map( G => n17728
                           , D => n13181, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_23_2_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_21_2_inst : DLH_X1 port map( G => n17726
                           , D => n13181, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_21_2_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_19_2_inst : DLH_X1 port map( G => n17724
                           , D => n13181, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_19_2_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_17_2_inst : DLH_X1 port map( G => n17722
                           , D => n13181, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_17_2_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_15_2_inst : DLH_X1 port map( G => n17720
                           , D => n13181, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_15_2_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_13_2_inst : DLH_X1 port map( G => n17718
                           , D => n13181, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_13_2_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_11_2_inst : DLH_X1 port map( G => n17716
                           , D => n13181, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_11_2_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_9_2_inst : DLH_X1 port map( G => n17714,
                           D => n13181, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_9_2_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_7_2_inst : DLH_X1 port map( G => n17712,
                           D => n13181, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_7_2_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_5_2_inst : DLH_X1 port map( G => n17710,
                           D => n13181, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_5_2_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_3_2_inst : DLH_X1 port map( G => n17708,
                           D => n13181, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_3_2_port);
   pipeline_RegFile_DEC_WB_RegBank_reg_1_2_inst : DLH_X1 port map( G => n17706,
                           D => n13181, Q => 
                           pipeline_RegFile_DEC_WB_RegBank_1_2_port);
   pipeline_IDEX_Stage_Reg2_out_IDEX_reg_2_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N136, CK => Clk, Q => n13811, QN
                           => n17497);
   pipeline_stageF_PC_reg_PC_out_reg_2_inst : DFFR_X1 port map( D => n3860, CK 
                           => Clk, RN => n17705, Q => n13810, QN => n7649);
   pipeline_IDEX_Stage_Reg1_out_IDEX_reg_2_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N104, CK => Clk, Q => n13809, QN
                           => net214731);
   pipeline_EXMEM_stage_DataToMem_out_EXMEM_reg_2_inst : DFF_X1 port map( D => 
                           pipeline_EXMEM_stage_N41, CK => Clk, Q => n13808, QN
                           => net214730);
   DataMem_Mem_reg_7_2_inst : DLH_X1 port map( G => n13079, D => DataMem_N2101,
                           Q => DataMem_Mem_7_2_port);
   DataMem_Mem_reg_6_2_inst : DLH_X1 port map( G => n13076, D => DataMem_N2037,
                           Q => DataMem_Mem_6_2_port);
   DataMem_Mem_reg_5_2_inst : DLH_X1 port map( G => n13073, D => DataMem_N1973,
                           Q => DataMem_Mem_5_2_port);
   DataMem_Mem_reg_4_2_inst : DLH_X1 port map( G => n13070, D => DataMem_N1909,
                           Q => DataMem_Mem_4_2_port);
   DataMem_Mem_reg_3_2_inst : DLH_X1 port map( G => n13067, D => DataMem_N1845,
                           Q => DataMem_Mem_3_2_port);
   DataMem_Mem_reg_2_2_inst : DLH_X1 port map( G => n13064, D => DataMem_N1781,
                           Q => DataMem_Mem_2_2_port);
   DataMem_Mem_reg_1_2_inst : DLH_X1 port map( G => n13061, D => DataMem_N1717,
                           Q => DataMem_Mem_1_2_port);
   DataMem_Mem_reg_0_2_inst : DLH_X1 port map( G => n13058, D => DataMem_N1653,
                           Q => DataMem_Mem_0_2_port);
   DataMem_Dataout_reg_2_inst : DLL_X1 port map( D => DataMem_N2167, GN => 
                           n17098, Q => DataMem_N2343);
   pipeline_EXMEM_stage_DataToMem_out_EXMEM_reg_3_inst : DFF_X1 port map( D => 
                           pipeline_EXMEM_stage_N42, CK => Clk, Q => n13807, QN
                           => net214729);
   DataMem_Mem_reg_7_3_inst : DLH_X1 port map( G => n13079, D => DataMem_N2103,
                           Q => DataMem_Mem_7_3_port);
   DataMem_Mem_reg_6_3_inst : DLH_X1 port map( G => n13076, D => DataMem_N2039,
                           Q => DataMem_Mem_6_3_port);
   DataMem_Mem_reg_5_3_inst : DLH_X1 port map( G => n13073, D => DataMem_N1975,
                           Q => DataMem_Mem_5_3_port);
   DataMem_Mem_reg_4_3_inst : DLH_X1 port map( G => n13070, D => DataMem_N1911,
                           Q => DataMem_Mem_4_3_port);
   DataMem_Mem_reg_3_3_inst : DLH_X1 port map( G => n13067, D => DataMem_N1847,
                           Q => DataMem_Mem_3_3_port);
   DataMem_Mem_reg_2_3_inst : DLH_X1 port map( G => n13064, D => DataMem_N1783,
                           Q => DataMem_Mem_2_3_port);
   DataMem_Mem_reg_1_3_inst : DLH_X1 port map( G => n13061, D => DataMem_N1719,
                           Q => DataMem_Mem_1_3_port);
   DataMem_Mem_reg_0_3_inst : DLH_X1 port map( G => n13058, D => DataMem_N1655,
                           Q => DataMem_Mem_0_3_port);
   DataMem_Dataout_reg_3_inst : DLL_X1 port map( D => DataMem_N2170, GN => 
                           n17098, Q => DataMem_N2340);
   pipeline_stageF_PC_reg_PC_out_reg_1_inst : DFFR_X1 port map( D => n3858, CK 
                           => Clk, RN => n17705, Q => n13806, QN => n7648);
   pipeline_EXMEM_stage_DataToMem_out_EXMEM_reg_1_inst : DFF_X1 port map( D => 
                           pipeline_EXMEM_stage_N40, CK => Clk, Q => n13805, QN
                           => net214728);
   pipeline_IDEX_Stage_Reg1_out_IDEX_reg_16_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N118, CK => Clk, Q => n13804, QN
                           => net214727);
   pipeline_EXMEM_stage_DataToMem_out_EXMEM_reg_16_inst : DFF_X1 port map( D =>
                           pipeline_EXMEM_stage_N55, CK => Clk, Q => n13803, QN
                           => net214726);
   DataMem_Mem_reg_7_16_inst : DLH_X1 port map( G => n13079, D => DataMem_N2129
                           , Q => DataMem_Mem_7_16_port);
   DataMem_Mem_reg_6_16_inst : DLH_X1 port map( G => n13076, D => DataMem_N2065
                           , Q => DataMem_Mem_6_16_port);
   DataMem_Mem_reg_5_16_inst : DLH_X1 port map( G => n13073, D => DataMem_N2001
                           , Q => DataMem_Mem_5_16_port);
   DataMem_Mem_reg_4_16_inst : DLH_X1 port map( G => n13070, D => DataMem_N1937
                           , Q => DataMem_Mem_4_16_port);
   DataMem_Mem_reg_3_16_inst : DLH_X1 port map( G => n13067, D => DataMem_N1873
                           , Q => DataMem_Mem_3_16_port);
   DataMem_Mem_reg_2_16_inst : DLH_X1 port map( G => n13064, D => DataMem_N1809
                           , Q => DataMem_Mem_2_16_port);
   DataMem_Mem_reg_1_16_inst : DLH_X1 port map( G => n13061, D => DataMem_N1745
                           , Q => DataMem_Mem_1_16_port);
   DataMem_Mem_reg_0_16_inst : DLH_X1 port map( G => n13058, D => DataMem_N1681
                           , Q => DataMem_Mem_0_16_port);
   DataMem_Dataout_reg_16_inst : DLL_X1 port map( D => DataMem_N2209, GN => 
                           n13055, Q => DataMem_N2301);
   pipeline_EXMEM_stage_DataToMem_out_EXMEM_reg_17_inst : DFF_X1 port map( D =>
                           pipeline_EXMEM_stage_N56, CK => Clk, Q => n13802, QN
                           => net214725);
   DataMem_Mem_reg_7_17_inst : DLH_X1 port map( G => n13079, D => DataMem_N2131
                           , Q => DataMem_Mem_7_17_port);
   DataMem_Mem_reg_6_17_inst : DLH_X1 port map( G => n13076, D => DataMem_N2067
                           , Q => DataMem_Mem_6_17_port);
   DataMem_Mem_reg_5_17_inst : DLH_X1 port map( G => n13073, D => DataMem_N2003
                           , Q => DataMem_Mem_5_17_port);
   DataMem_Mem_reg_4_17_inst : DLH_X1 port map( G => n13070, D => DataMem_N1939
                           , Q => DataMem_Mem_4_17_port);
   DataMem_Mem_reg_3_17_inst : DLH_X1 port map( G => n13067, D => DataMem_N1875
                           , Q => DataMem_Mem_3_17_port);
   DataMem_Mem_reg_2_17_inst : DLH_X1 port map( G => n13064, D => DataMem_N1811
                           , Q => DataMem_Mem_2_17_port);
   DataMem_Mem_reg_1_17_inst : DLH_X1 port map( G => n13061, D => DataMem_N1747
                           , Q => DataMem_Mem_1_17_port);
   DataMem_Mem_reg_0_17_inst : DLH_X1 port map( G => n13058, D => DataMem_N1683
                           , Q => DataMem_Mem_0_17_port);
   DataMem_Dataout_reg_17_inst : DLL_X1 port map( D => DataMem_N2212, GN => 
                           n13055, Q => DataMem_N2298);
   pipeline_EXMEM_stage_DataToMem_out_EXMEM_reg_18_inst : DFF_X1 port map( D =>
                           pipeline_EXMEM_stage_N57, CK => Clk, Q => n13801, QN
                           => net214724);
   DataMem_Mem_reg_7_18_inst : DLH_X1 port map( G => n13079, D => DataMem_N2133
                           , Q => DataMem_Mem_7_18_port);
   DataMem_Mem_reg_6_18_inst : DLH_X1 port map( G => n13076, D => DataMem_N2069
                           , Q => DataMem_Mem_6_18_port);
   DataMem_Mem_reg_5_18_inst : DLH_X1 port map( G => n13073, D => DataMem_N2005
                           , Q => DataMem_Mem_5_18_port);
   DataMem_Mem_reg_4_18_inst : DLH_X1 port map( G => n13070, D => DataMem_N1941
                           , Q => DataMem_Mem_4_18_port);
   DataMem_Mem_reg_3_18_inst : DLH_X1 port map( G => n13067, D => DataMem_N1877
                           , Q => DataMem_Mem_3_18_port);
   DataMem_Mem_reg_2_18_inst : DLH_X1 port map( G => n13064, D => DataMem_N1813
                           , Q => DataMem_Mem_2_18_port);
   DataMem_Mem_reg_1_18_inst : DLH_X1 port map( G => n13061, D => DataMem_N1749
                           , Q => DataMem_Mem_1_18_port);
   DataMem_Mem_reg_0_18_inst : DLH_X1 port map( G => n13058, D => DataMem_N1685
                           , Q => DataMem_Mem_0_18_port);
   DataMem_Dataout_reg_18_inst : DLL_X1 port map( D => DataMem_N2215, GN => 
                           n17098, Q => DataMem_N2295);
   pipeline_EXMEM_stage_DataToMem_out_EXMEM_reg_19_inst : DFF_X1 port map( D =>
                           pipeline_EXMEM_stage_N58, CK => Clk, Q => n13800, QN
                           => net214723);
   DataMem_Mem_reg_7_19_inst : DLH_X1 port map( G => n13079, D => DataMem_N2135
                           , Q => DataMem_Mem_7_19_port);
   DataMem_Mem_reg_6_19_inst : DLH_X1 port map( G => n13076, D => DataMem_N2071
                           , Q => DataMem_Mem_6_19_port);
   DataMem_Mem_reg_5_19_inst : DLH_X1 port map( G => n13073, D => DataMem_N2007
                           , Q => DataMem_Mem_5_19_port);
   DataMem_Mem_reg_4_19_inst : DLH_X1 port map( G => n13070, D => DataMem_N1943
                           , Q => DataMem_Mem_4_19_port);
   DataMem_Mem_reg_3_19_inst : DLH_X1 port map( G => n13067, D => DataMem_N1879
                           , Q => DataMem_Mem_3_19_port);
   DataMem_Mem_reg_2_19_inst : DLH_X1 port map( G => n13064, D => DataMem_N1815
                           , Q => DataMem_Mem_2_19_port);
   DataMem_Mem_reg_1_19_inst : DLH_X1 port map( G => n13061, D => DataMem_N1751
                           , Q => DataMem_Mem_1_19_port);
   DataMem_Mem_reg_0_19_inst : DLH_X1 port map( G => n13058, D => DataMem_N1687
                           , Q => DataMem_Mem_0_19_port);
   DataMem_Dataout_reg_19_inst : DLL_X1 port map( D => DataMem_N2218, GN => 
                           n13055, Q => DataMem_N2292);
   pipeline_EXMEM_stage_DataToMem_out_EXMEM_reg_20_inst : DFF_X1 port map( D =>
                           pipeline_EXMEM_stage_N59, CK => Clk, Q => n13799, QN
                           => net214722);
   DataMem_Mem_reg_7_20_inst : DLH_X1 port map( G => n13079, D => DataMem_N2137
                           , Q => DataMem_Mem_7_20_port);
   DataMem_Mem_reg_6_20_inst : DLH_X1 port map( G => n13076, D => DataMem_N2073
                           , Q => DataMem_Mem_6_20_port);
   DataMem_Mem_reg_5_20_inst : DLH_X1 port map( G => n13073, D => DataMem_N2009
                           , Q => DataMem_Mem_5_20_port);
   DataMem_Mem_reg_4_20_inst : DLH_X1 port map( G => n13070, D => DataMem_N1945
                           , Q => DataMem_Mem_4_20_port);
   DataMem_Mem_reg_3_20_inst : DLH_X1 port map( G => n13067, D => DataMem_N1881
                           , Q => DataMem_Mem_3_20_port);
   DataMem_Mem_reg_2_20_inst : DLH_X1 port map( G => n13064, D => DataMem_N1817
                           , Q => DataMem_Mem_2_20_port);
   DataMem_Mem_reg_1_20_inst : DLH_X1 port map( G => n13061, D => DataMem_N1753
                           , Q => DataMem_Mem_1_20_port);
   DataMem_Mem_reg_0_20_inst : DLH_X1 port map( G => n13058, D => DataMem_N1689
                           , Q => DataMem_Mem_0_20_port);
   DataMem_Dataout_reg_20_inst : DLL_X1 port map( D => DataMem_N2221, GN => 
                           n17098, Q => DataMem_N2289);
   pipeline_EXMEM_stage_DataToMem_out_EXMEM_reg_21_inst : DFF_X1 port map( D =>
                           pipeline_EXMEM_stage_N60, CK => Clk, Q => n13798, QN
                           => net214721);
   DataMem_Mem_reg_7_21_inst : DLH_X1 port map( G => n13079, D => DataMem_N2139
                           , Q => DataMem_Mem_7_21_port);
   DataMem_Mem_reg_6_21_inst : DLH_X1 port map( G => n13076, D => DataMem_N2075
                           , Q => DataMem_Mem_6_21_port);
   DataMem_Mem_reg_5_21_inst : DLH_X1 port map( G => n13073, D => DataMem_N2011
                           , Q => DataMem_Mem_5_21_port);
   DataMem_Mem_reg_4_21_inst : DLH_X1 port map( G => n13070, D => DataMem_N1947
                           , Q => DataMem_Mem_4_21_port);
   DataMem_Mem_reg_3_21_inst : DLH_X1 port map( G => n13067, D => DataMem_N1883
                           , Q => DataMem_Mem_3_21_port);
   DataMem_Mem_reg_2_21_inst : DLH_X1 port map( G => n13064, D => DataMem_N1819
                           , Q => DataMem_Mem_2_21_port);
   DataMem_Mem_reg_1_21_inst : DLH_X1 port map( G => n13061, D => DataMem_N1755
                           , Q => DataMem_Mem_1_21_port);
   DataMem_Mem_reg_0_21_inst : DLH_X1 port map( G => n13058, D => DataMem_N1691
                           , Q => DataMem_Mem_0_21_port);
   DataMem_Dataout_reg_21_inst : DLL_X1 port map( D => DataMem_N2224, GN => 
                           n17098, Q => DataMem_N2286);
   pipeline_EXMEM_stage_DataToMem_out_EXMEM_reg_22_inst : DFF_X1 port map( D =>
                           pipeline_EXMEM_stage_N61, CK => Clk, Q => n13797, QN
                           => net214720);
   DataMem_Mem_reg_7_22_inst : DLH_X1 port map( G => n13079, D => DataMem_N2141
                           , Q => DataMem_Mem_7_22_port);
   DataMem_Mem_reg_6_22_inst : DLH_X1 port map( G => n13076, D => DataMem_N2077
                           , Q => DataMem_Mem_6_22_port);
   DataMem_Mem_reg_5_22_inst : DLH_X1 port map( G => n13073, D => DataMem_N2013
                           , Q => DataMem_Mem_5_22_port);
   DataMem_Mem_reg_4_22_inst : DLH_X1 port map( G => n13070, D => DataMem_N1949
                           , Q => DataMem_Mem_4_22_port);
   DataMem_Mem_reg_3_22_inst : DLH_X1 port map( G => n13067, D => DataMem_N1885
                           , Q => DataMem_Mem_3_22_port);
   DataMem_Mem_reg_2_22_inst : DLH_X1 port map( G => n13064, D => DataMem_N1821
                           , Q => DataMem_Mem_2_22_port);
   DataMem_Mem_reg_1_22_inst : DLH_X1 port map( G => n13061, D => DataMem_N1757
                           , Q => DataMem_Mem_1_22_port);
   DataMem_Mem_reg_0_22_inst : DLH_X1 port map( G => n13058, D => DataMem_N1693
                           , Q => DataMem_Mem_0_22_port);
   DataMem_Dataout_reg_22_inst : DLL_X1 port map( D => DataMem_N2227, GN => 
                           n13055, Q => DataMem_N2283);
   pipeline_EXMEM_stage_DataToMem_out_EXMEM_reg_23_inst : DFF_X1 port map( D =>
                           pipeline_EXMEM_stage_N62, CK => Clk, Q => n13796, QN
                           => net214719);
   DataMem_Mem_reg_7_23_inst : DLH_X1 port map( G => n13079, D => DataMem_N2143
                           , Q => DataMem_Mem_7_23_port);
   DataMem_Mem_reg_6_23_inst : DLH_X1 port map( G => n13076, D => DataMem_N2079
                           , Q => DataMem_Mem_6_23_port);
   DataMem_Mem_reg_5_23_inst : DLH_X1 port map( G => n13073, D => DataMem_N2015
                           , Q => DataMem_Mem_5_23_port);
   DataMem_Mem_reg_4_23_inst : DLH_X1 port map( G => n13070, D => DataMem_N1951
                           , Q => DataMem_Mem_4_23_port);
   DataMem_Mem_reg_3_23_inst : DLH_X1 port map( G => n13067, D => DataMem_N1887
                           , Q => DataMem_Mem_3_23_port);
   DataMem_Mem_reg_2_23_inst : DLH_X1 port map( G => n13064, D => DataMem_N1823
                           , Q => DataMem_Mem_2_23_port);
   DataMem_Mem_reg_1_23_inst : DLH_X1 port map( G => n13061, D => DataMem_N1759
                           , Q => DataMem_Mem_1_23_port);
   DataMem_Mem_reg_0_23_inst : DLH_X1 port map( G => n13058, D => DataMem_N1695
                           , Q => DataMem_Mem_0_23_port);
   DataMem_Dataout_reg_23_inst : DLL_X1 port map( D => DataMem_N2230, GN => 
                           n13055, Q => DataMem_N2280);
   pipeline_EXMEM_stage_DataToMem_out_EXMEM_reg_25_inst : DFF_X1 port map( D =>
                           pipeline_EXMEM_stage_N64, CK => Clk, Q => n13795, QN
                           => net214718);
   DataMem_Mem_reg_7_25_inst : DLH_X1 port map( G => n13079, D => DataMem_N2147
                           , Q => DataMem_Mem_7_25_port);
   DataMem_Mem_reg_6_25_inst : DLH_X1 port map( G => n13076, D => DataMem_N2083
                           , Q => DataMem_Mem_6_25_port);
   DataMem_Mem_reg_5_25_inst : DLH_X1 port map( G => n13073, D => DataMem_N2019
                           , Q => DataMem_Mem_5_25_port);
   DataMem_Mem_reg_4_25_inst : DLH_X1 port map( G => n13070, D => DataMem_N1955
                           , Q => DataMem_Mem_4_25_port);
   DataMem_Mem_reg_3_25_inst : DLH_X1 port map( G => n13067, D => DataMem_N1891
                           , Q => DataMem_Mem_3_25_port);
   DataMem_Mem_reg_2_25_inst : DLH_X1 port map( G => n13064, D => DataMem_N1827
                           , Q => DataMem_Mem_2_25_port);
   DataMem_Mem_reg_1_25_inst : DLH_X1 port map( G => n13061, D => DataMem_N1763
                           , Q => DataMem_Mem_1_25_port);
   DataMem_Mem_reg_0_25_inst : DLH_X1 port map( G => n13058, D => DataMem_N1699
                           , Q => DataMem_Mem_0_25_port);
   DataMem_Dataout_reg_25_inst : DLL_X1 port map( D => DataMem_N2236, GN => 
                           n17098, Q => DataMem_N2274);
   pipeline_EXMEM_stage_DataToMem_out_EXMEM_reg_26_inst : DFF_X1 port map( D =>
                           pipeline_EXMEM_stage_N65, CK => Clk, Q => n13794, QN
                           => net214717);
   DataMem_Mem_reg_7_26_inst : DLH_X1 port map( G => n13079, D => DataMem_N2149
                           , Q => DataMem_Mem_7_26_port);
   DataMem_Mem_reg_6_26_inst : DLH_X1 port map( G => n13076, D => DataMem_N2085
                           , Q => DataMem_Mem_6_26_port);
   DataMem_Mem_reg_5_26_inst : DLH_X1 port map( G => n13073, D => DataMem_N2021
                           , Q => DataMem_Mem_5_26_port);
   DataMem_Mem_reg_4_26_inst : DLH_X1 port map( G => n13070, D => DataMem_N1957
                           , Q => DataMem_Mem_4_26_port);
   DataMem_Mem_reg_3_26_inst : DLH_X1 port map( G => n13067, D => DataMem_N1893
                           , Q => DataMem_Mem_3_26_port);
   DataMem_Mem_reg_2_26_inst : DLH_X1 port map( G => n13064, D => DataMem_N1829
                           , Q => DataMem_Mem_2_26_port);
   DataMem_Mem_reg_1_26_inst : DLH_X1 port map( G => n13061, D => DataMem_N1765
                           , Q => DataMem_Mem_1_26_port);
   DataMem_Mem_reg_0_26_inst : DLH_X1 port map( G => n13058, D => DataMem_N1701
                           , Q => DataMem_Mem_0_26_port);
   DataMem_Dataout_reg_26_inst : DLL_X1 port map( D => DataMem_N2239, GN => 
                           n17098, Q => DataMem_N2271);
   pipeline_EXMEM_stage_DataToMem_out_EXMEM_reg_27_inst : DFF_X1 port map( D =>
                           pipeline_EXMEM_stage_N66, CK => Clk, Q => n13793, QN
                           => net214716);
   DataMem_Mem_reg_7_27_inst : DLH_X1 port map( G => n13079, D => DataMem_N2151
                           , Q => DataMem_Mem_7_27_port);
   DataMem_Mem_reg_6_27_inst : DLH_X1 port map( G => n13076, D => DataMem_N2087
                           , Q => DataMem_Mem_6_27_port);
   DataMem_Mem_reg_5_27_inst : DLH_X1 port map( G => n13073, D => DataMem_N2023
                           , Q => DataMem_Mem_5_27_port);
   DataMem_Mem_reg_4_27_inst : DLH_X1 port map( G => n13070, D => DataMem_N1959
                           , Q => DataMem_Mem_4_27_port);
   DataMem_Mem_reg_3_27_inst : DLH_X1 port map( G => n13067, D => DataMem_N1895
                           , Q => DataMem_Mem_3_27_port);
   DataMem_Mem_reg_2_27_inst : DLH_X1 port map( G => n13064, D => DataMem_N1831
                           , Q => DataMem_Mem_2_27_port);
   DataMem_Mem_reg_1_27_inst : DLH_X1 port map( G => n13061, D => DataMem_N1767
                           , Q => DataMem_Mem_1_27_port);
   DataMem_Mem_reg_0_27_inst : DLH_X1 port map( G => n13058, D => DataMem_N1703
                           , Q => DataMem_Mem_0_27_port);
   DataMem_Dataout_reg_27_inst : DLL_X1 port map( D => DataMem_N2242, GN => 
                           n17098, Q => DataMem_N2268);
   pipeline_EXMEM_stage_DataToMem_out_EXMEM_reg_29_inst : DFF_X1 port map( D =>
                           pipeline_EXMEM_stage_N68, CK => Clk, Q => n13792, QN
                           => net214715);
   DataMem_Mem_reg_7_29_inst : DLH_X1 port map( G => n13079, D => DataMem_N2155
                           , Q => DataMem_Mem_7_29_port);
   DataMem_Mem_reg_6_29_inst : DLH_X1 port map( G => n13076, D => DataMem_N2091
                           , Q => DataMem_Mem_6_29_port);
   DataMem_Mem_reg_5_29_inst : DLH_X1 port map( G => n13073, D => DataMem_N2027
                           , Q => DataMem_Mem_5_29_port);
   DataMem_Mem_reg_4_29_inst : DLH_X1 port map( G => n13070, D => DataMem_N1963
                           , Q => DataMem_Mem_4_29_port);
   DataMem_Mem_reg_3_29_inst : DLH_X1 port map( G => n13067, D => DataMem_N1899
                           , Q => DataMem_Mem_3_29_port);
   DataMem_Mem_reg_2_29_inst : DLH_X1 port map( G => n13064, D => DataMem_N1835
                           , Q => DataMem_Mem_2_29_port);
   DataMem_Mem_reg_1_29_inst : DLH_X1 port map( G => n13061, D => DataMem_N1771
                           , Q => DataMem_Mem_1_29_port);
   DataMem_Mem_reg_0_29_inst : DLH_X1 port map( G => n13058, D => DataMem_N1707
                           , Q => DataMem_Mem_0_29_port);
   DataMem_Dataout_reg_29_inst : DLL_X1 port map( D => DataMem_N2248, GN => 
                           n17098, Q => DataMem_N2262);
   pipeline_EXMEM_stage_DataToMem_out_EXMEM_reg_30_inst : DFF_X1 port map( D =>
                           pipeline_EXMEM_stage_N69, CK => Clk, Q => n13791, QN
                           => net214714);
   DataMem_Mem_reg_7_30_inst : DLH_X1 port map( G => n13079, D => DataMem_N2157
                           , Q => DataMem_Mem_7_30_port);
   DataMem_Mem_reg_6_30_inst : DLH_X1 port map( G => n13076, D => DataMem_N2093
                           , Q => DataMem_Mem_6_30_port);
   DataMem_Mem_reg_5_30_inst : DLH_X1 port map( G => n13073, D => DataMem_N2029
                           , Q => DataMem_Mem_5_30_port);
   DataMem_Mem_reg_4_30_inst : DLH_X1 port map( G => n13070, D => DataMem_N1965
                           , Q => DataMem_Mem_4_30_port);
   DataMem_Mem_reg_3_30_inst : DLH_X1 port map( G => n13067, D => DataMem_N1901
                           , Q => DataMem_Mem_3_30_port);
   DataMem_Mem_reg_2_30_inst : DLH_X1 port map( G => n13064, D => DataMem_N1837
                           , Q => DataMem_Mem_2_30_port);
   DataMem_Mem_reg_1_30_inst : DLH_X1 port map( G => n13061, D => DataMem_N1773
                           , Q => DataMem_Mem_1_30_port);
   DataMem_Mem_reg_0_30_inst : DLH_X1 port map( G => n13058, D => DataMem_N1709
                           , Q => DataMem_Mem_0_30_port);
   DataMem_Dataout_reg_30_inst : DLL_X1 port map( D => DataMem_N2251, GN => 
                           n17098, Q => DataMem_N2259);
   pipeline_EXMEM_stage_DataToMem_out_EXMEM_reg_13_inst : DFF_X1 port map( D =>
                           pipeline_EXMEM_stage_N52, CK => Clk, Q => n13790, QN
                           => net214713);
   DataMem_Mem_reg_7_13_inst : DLH_X1 port map( G => n13079, D => DataMem_N2123
                           , Q => DataMem_Mem_7_13_port);
   DataMem_Mem_reg_6_13_inst : DLH_X1 port map( G => n13076, D => DataMem_N2059
                           , Q => DataMem_Mem_6_13_port);
   DataMem_Mem_reg_5_13_inst : DLH_X1 port map( G => n13073, D => DataMem_N1995
                           , Q => DataMem_Mem_5_13_port);
   DataMem_Mem_reg_4_13_inst : DLH_X1 port map( G => n13070, D => DataMem_N1931
                           , Q => DataMem_Mem_4_13_port);
   DataMem_Mem_reg_3_13_inst : DLH_X1 port map( G => n13067, D => DataMem_N1867
                           , Q => DataMem_Mem_3_13_port);
   DataMem_Mem_reg_2_13_inst : DLH_X1 port map( G => n13064, D => DataMem_N1803
                           , Q => DataMem_Mem_2_13_port);
   DataMem_Mem_reg_1_13_inst : DLH_X1 port map( G => n13061, D => DataMem_N1739
                           , Q => DataMem_Mem_1_13_port);
   DataMem_Mem_reg_0_13_inst : DLH_X1 port map( G => n13058, D => DataMem_N1675
                           , Q => DataMem_Mem_0_13_port);
   DataMem_Dataout_reg_13_inst : DLL_X1 port map( D => DataMem_N2200, GN => 
                           n13055, Q => DataMem_N2310);
   pipeline_EXMEM_stage_DataToMem_out_EXMEM_reg_15_inst : DFF_X1 port map( D =>
                           pipeline_EXMEM_stage_N54, CK => Clk, Q => n13789, QN
                           => net214712);
   DataMem_Mem_reg_7_15_inst : DLH_X1 port map( G => n13079, D => DataMem_N2127
                           , Q => DataMem_Mem_7_15_port);
   DataMem_Mem_reg_6_15_inst : DLH_X1 port map( G => n13076, D => DataMem_N2063
                           , Q => DataMem_Mem_6_15_port);
   DataMem_Mem_reg_5_15_inst : DLH_X1 port map( G => n13073, D => DataMem_N1999
                           , Q => DataMem_Mem_5_15_port);
   DataMem_Mem_reg_4_15_inst : DLH_X1 port map( G => n13070, D => DataMem_N1935
                           , Q => DataMem_Mem_4_15_port);
   DataMem_Mem_reg_3_15_inst : DLH_X1 port map( G => n13067, D => DataMem_N1871
                           , Q => DataMem_Mem_3_15_port);
   DataMem_Mem_reg_2_15_inst : DLH_X1 port map( G => n13064, D => DataMem_N1807
                           , Q => DataMem_Mem_2_15_port);
   DataMem_Mem_reg_1_15_inst : DLH_X1 port map( G => n13061, D => DataMem_N1743
                           , Q => DataMem_Mem_1_15_port);
   DataMem_Mem_reg_0_15_inst : DLH_X1 port map( G => n13058, D => DataMem_N1679
                           , Q => DataMem_Mem_0_15_port);
   DataMem_Dataout_reg_15_inst : DLL_X1 port map( D => DataMem_N2206, GN => 
                           n13055, Q => DataMem_N2304);
   pipeline_EXMEM_stage_DataToMem_out_EXMEM_reg_14_inst : DFF_X1 port map( D =>
                           pipeline_EXMEM_stage_N53, CK => Clk, Q => n13788, QN
                           => net214711);
   DataMem_Mem_reg_7_14_inst : DLH_X1 port map( G => n13079, D => DataMem_N2125
                           , Q => DataMem_Mem_7_14_port);
   DataMem_Mem_reg_6_14_inst : DLH_X1 port map( G => n13076, D => DataMem_N2061
                           , Q => DataMem_Mem_6_14_port);
   DataMem_Mem_reg_5_14_inst : DLH_X1 port map( G => n13073, D => DataMem_N1997
                           , Q => DataMem_Mem_5_14_port);
   DataMem_Mem_reg_4_14_inst : DLH_X1 port map( G => n13070, D => DataMem_N1933
                           , Q => DataMem_Mem_4_14_port);
   DataMem_Mem_reg_3_14_inst : DLH_X1 port map( G => n13067, D => DataMem_N1869
                           , Q => DataMem_Mem_3_14_port);
   DataMem_Mem_reg_2_14_inst : DLH_X1 port map( G => n13064, D => DataMem_N1805
                           , Q => DataMem_Mem_2_14_port);
   DataMem_Mem_reg_1_14_inst : DLH_X1 port map( G => n13061, D => DataMem_N1741
                           , Q => DataMem_Mem_1_14_port);
   DataMem_Mem_reg_0_14_inst : DLH_X1 port map( G => n13058, D => DataMem_N1677
                           , Q => DataMem_Mem_0_14_port);
   DataMem_Dataout_reg_14_inst : DLL_X1 port map( D => DataMem_N2203, GN => 
                           n13055, Q => DataMem_N2307);
   pipeline_EXMEM_stage_DataToMem_out_EXMEM_reg_28_inst : DFF_X1 port map( D =>
                           pipeline_EXMEM_stage_N67, CK => Clk, Q => n13787, QN
                           => net214710);
   DataMem_Mem_reg_7_28_inst : DLH_X1 port map( G => n13079, D => DataMem_N2153
                           , Q => DataMem_Mem_7_28_port);
   DataMem_Mem_reg_6_28_inst : DLH_X1 port map( G => n13076, D => DataMem_N2089
                           , Q => DataMem_Mem_6_28_port);
   DataMem_Mem_reg_5_28_inst : DLH_X1 port map( G => n13073, D => DataMem_N2025
                           , Q => DataMem_Mem_5_28_port);
   DataMem_Mem_reg_4_28_inst : DLH_X1 port map( G => n13070, D => DataMem_N1961
                           , Q => DataMem_Mem_4_28_port);
   DataMem_Mem_reg_3_28_inst : DLH_X1 port map( G => n13067, D => DataMem_N1897
                           , Q => DataMem_Mem_3_28_port);
   DataMem_Mem_reg_2_28_inst : DLH_X1 port map( G => n13064, D => DataMem_N1833
                           , Q => DataMem_Mem_2_28_port);
   DataMem_Mem_reg_1_28_inst : DLH_X1 port map( G => n13061, D => DataMem_N1769
                           , Q => DataMem_Mem_1_28_port);
   DataMem_Mem_reg_0_28_inst : DLH_X1 port map( G => n13058, D => DataMem_N1705
                           , Q => DataMem_Mem_0_28_port);
   DataMem_Dataout_reg_28_inst : DLL_X1 port map( D => DataMem_N2245, GN => 
                           n17098, Q => DataMem_N2265);
   pipeline_EXMEM_stage_DataToMem_out_EXMEM_reg_24_inst : DFF_X1 port map( D =>
                           pipeline_EXMEM_stage_N63, CK => Clk, Q => n13786, QN
                           => net214709);
   DataMem_Mem_reg_7_24_inst : DLH_X1 port map( G => n13079, D => DataMem_N2145
                           , Q => DataMem_Mem_7_24_port);
   DataMem_Mem_reg_6_24_inst : DLH_X1 port map( G => n13076, D => DataMem_N2081
                           , Q => DataMem_Mem_6_24_port);
   DataMem_Mem_reg_5_24_inst : DLH_X1 port map( G => n13073, D => DataMem_N2017
                           , Q => DataMem_Mem_5_24_port);
   DataMem_Mem_reg_4_24_inst : DLH_X1 port map( G => n13070, D => DataMem_N1953
                           , Q => DataMem_Mem_4_24_port);
   DataMem_Mem_reg_3_24_inst : DLH_X1 port map( G => n13067, D => DataMem_N1889
                           , Q => DataMem_Mem_3_24_port);
   DataMem_Mem_reg_2_24_inst : DLH_X1 port map( G => n13064, D => DataMem_N1825
                           , Q => DataMem_Mem_2_24_port);
   DataMem_Mem_reg_1_24_inst : DLH_X1 port map( G => n13061, D => DataMem_N1761
                           , Q => DataMem_Mem_1_24_port);
   DataMem_Mem_reg_0_24_inst : DLH_X1 port map( G => n13058, D => DataMem_N1697
                           , Q => DataMem_Mem_0_24_port);
   DataMem_Dataout_reg_24_inst : DLL_X1 port map( D => DataMem_N2233, GN => 
                           n13055, Q => DataMem_N2277);
   pipeline_EXMEM_stage_DataToMem_out_EXMEM_reg_8_inst : DFF_X1 port map( D => 
                           pipeline_EXMEM_stage_N47, CK => Clk, Q => n13785, QN
                           => net214708);
   DataMem_Mem_reg_7_8_inst : DLH_X1 port map( G => n13079, D => DataMem_N2113,
                           Q => DataMem_Mem_7_8_port);
   DataMem_Mem_reg_6_8_inst : DLH_X1 port map( G => n13076, D => DataMem_N2049,
                           Q => DataMem_Mem_6_8_port);
   DataMem_Mem_reg_5_8_inst : DLH_X1 port map( G => n13073, D => DataMem_N1985,
                           Q => DataMem_Mem_5_8_port);
   DataMem_Mem_reg_4_8_inst : DLH_X1 port map( G => n13070, D => DataMem_N1921,
                           Q => DataMem_Mem_4_8_port);
   DataMem_Mem_reg_3_8_inst : DLH_X1 port map( G => n13067, D => DataMem_N1857,
                           Q => DataMem_Mem_3_8_port);
   DataMem_Mem_reg_2_8_inst : DLH_X1 port map( G => n13064, D => DataMem_N1793,
                           Q => DataMem_Mem_2_8_port);
   DataMem_Mem_reg_1_8_inst : DLH_X1 port map( G => n13061, D => DataMem_N1729,
                           Q => DataMem_Mem_1_8_port);
   DataMem_Mem_reg_0_8_inst : DLH_X1 port map( G => n13058, D => DataMem_N1665,
                           Q => DataMem_Mem_0_8_port);
   DataMem_Dataout_reg_8_inst : DLL_X1 port map( D => DataMem_N2185, GN => 
                           n17098, Q => DataMem_N2325);
   pipeline_EXMEM_stage_DataToMem_out_EXMEM_reg_0_inst : DFF_X1 port map( D => 
                           pipeline_EXMEM_stage_N39, CK => Clk, Q => n13784, QN
                           => net214707);
   DataMem_Mem_reg_7_0_inst : DLH_X1 port map( G => n13079, D => DataMem_N2097,
                           Q => DataMem_Mem_7_0_port);
   DataMem_Mem_reg_6_0_inst : DLH_X1 port map( G => n13076, D => DataMem_N2033,
                           Q => DataMem_Mem_6_0_port);
   DataMem_Mem_reg_5_0_inst : DLH_X1 port map( G => n13073, D => DataMem_N1969,
                           Q => DataMem_Mem_5_0_port);
   DataMem_Mem_reg_4_0_inst : DLH_X1 port map( G => n13070, D => DataMem_N1905,
                           Q => DataMem_Mem_4_0_port);
   DataMem_Mem_reg_3_0_inst : DLH_X1 port map( G => n13067, D => DataMem_N1841,
                           Q => DataMem_Mem_3_0_port);
   DataMem_Mem_reg_2_0_inst : DLH_X1 port map( G => n13064, D => DataMem_N1777,
                           Q => DataMem_Mem_2_0_port);
   DataMem_Mem_reg_1_0_inst : DLH_X1 port map( G => n13061, D => DataMem_N1713,
                           Q => DataMem_Mem_1_0_port);
   DataMem_Mem_reg_0_0_inst : DLH_X1 port map( G => n13058, D => DataMem_N1649,
                           Q => DataMem_Mem_0_0_port);
   DataMem_Dataout_reg_0_inst : DLL_X1 port map( D => DataMem_N2161, GN => 
                           n17098, Q => DataMem_N2349);
   pipeline_EXMEM_stage_DataToMem_out_EXMEM_reg_31_inst : DFF_X1 port map( D =>
                           pipeline_EXMEM_stage_N70, CK => Clk, Q => n13783, QN
                           => net214706);
   DataMem_Mem_reg_6_31_inst : DLH_X1 port map( G => n13076, D => DataMem_N2095
                           , Q => DataMem_Mem_6_31_port);
   DataMem_Mem_reg_5_31_inst : DLH_X1 port map( G => n13073, D => DataMem_N2031
                           , Q => DataMem_Mem_5_31_port);
   DataMem_Mem_reg_4_31_inst : DLH_X1 port map( G => n13070, D => DataMem_N1967
                           , Q => DataMem_Mem_4_31_port);
   DataMem_Mem_reg_3_31_inst : DLH_X1 port map( G => n13067, D => DataMem_N1903
                           , Q => DataMem_Mem_3_31_port);
   DataMem_Mem_reg_2_31_inst : DLH_X1 port map( G => n13064, D => DataMem_N1839
                           , Q => DataMem_Mem_2_31_port);
   DataMem_Mem_reg_1_31_inst : DLH_X1 port map( G => n13061, D => DataMem_N1775
                           , Q => DataMem_Mem_1_31_port);
   DataMem_Mem_reg_0_31_inst : DLH_X1 port map( G => n13058, D => DataMem_N1711
                           , Q => DataMem_Mem_0_31_port);
   n415 <= '0';
   pipeline_stageM_Addr_to_Dram_reg_4_inst : DLL_X1 port map( D => 
                           pipeline_Alu_Out_Addr_to_mem_4_port, GN => n12766, Q
                           => addr_to_dataRam_4_port);
   pipeline_IDEX_Stage_EXE_controls_out_IDEX_reg_1_inst : DFF_X2 port map( D =>
                           pipeline_IDEX_Stage_N94, CK => Clk, Q => 
                           pipeline_stageE_EXE_ALU_add_alu_sCout_0_port, QN => 
                           n17381);
   pipeline_stageM_Addr_to_Dram_reg_3_inst : DLL_X1 port map( D => 
                           pipeline_Alu_Out_Addr_to_mem_3_port, GN => n17155, Q
                           => addr_to_dataRam_3_port);
   pipeline_stageM_Addr_to_Dram_reg_2_inst : DLL_X1 port map( D => 
                           pipeline_Alu_Out_Addr_to_mem_2_port, GN => n12766, Q
                           => addr_to_dataRam_2_port);
   U4372 : TINV_X1 port map( I => n7676, EN => pipeline_stageF_PC_reg_N0, ZN =>
                           addr_to_iram_31_port);
   U4374 : TINV_X1 port map( I => n7649, EN => pipeline_stageF_PC_reg_N29, ZN 
                           => addr_to_iram_2_port);
   U4375 : TINV_X1 port map( I => n7659, EN => pipeline_stageF_PC_reg_N31, ZN 
                           => pipeline_stageF_PC_plus4_N7);
   U4376 : TINV_X1 port map( I => n7648, EN => pipeline_stageF_PC_reg_N30, ZN 
                           => pipeline_stageF_PC_plus4_N8);
   U4377 : TINV_X1 port map( I => n7658, EN => pipeline_stageF_PC_reg_N28, ZN 
                           => addr_to_iram_3_port);
   U4378 : TINV_X1 port map( I => n7656, EN => pipeline_stageF_PC_reg_N27, ZN 
                           => addr_to_iram_4_port);
   U4379 : TINV_X1 port map( I => n7655, EN => pipeline_stageF_PC_reg_N26, ZN 
                           => addr_to_iram_5_port);
   U4380 : TINV_X1 port map( I => n7654, EN => pipeline_stageF_PC_reg_N25, ZN 
                           => addr_to_iram_6_port);
   U4381 : TINV_X1 port map( I => n7657, EN => pipeline_stageF_PC_reg_N24, ZN 
                           => addr_to_iram_7_port);
   U4382 : TINV_X1 port map( I => n7660, EN => pipeline_stageF_PC_reg_N23, ZN 
                           => addr_to_iram_8_port);
   U4383 : TINV_X1 port map( I => n7652, EN => pipeline_stageF_PC_reg_N22, ZN 
                           => addr_to_iram_9_port);
   U4384 : TINV_X1 port map( I => n7651, EN => pipeline_stageF_PC_reg_N21, ZN 
                           => addr_to_iram_10_port);
   U4385 : TINV_X1 port map( I => n7653, EN => pipeline_stageF_PC_reg_N20, ZN 
                           => addr_to_iram_11_port);
   U4386 : TINV_X1 port map( I => n7650, EN => pipeline_stageF_PC_reg_N19, ZN 
                           => addr_to_iram_12_port);
   U4387 : TINV_X1 port map( I => n7661, EN => pipeline_stageF_PC_reg_N18, ZN 
                           => addr_to_iram_13_port);
   U4388 : TINV_X1 port map( I => n7662, EN => pipeline_stageF_PC_reg_N17, ZN 
                           => addr_to_iram_14_port);
   U4389 : TINV_X1 port map( I => n7663, EN => pipeline_stageF_PC_reg_N16, ZN 
                           => addr_to_iram_15_port);
   U4390 : TINV_X1 port map( I => n7711, EN => pipeline_stageF_PC_reg_N15, ZN 
                           => addr_to_iram_16_port);
   U4391 : TINV_X1 port map( I => n7664, EN => pipeline_stageF_PC_reg_N14, ZN 
                           => addr_to_iram_17_port);
   U4392 : TINV_X1 port map( I => n7665, EN => pipeline_stageF_PC_reg_N13, ZN 
                           => addr_to_iram_18_port);
   U4393 : TINV_X1 port map( I => n7666, EN => pipeline_stageF_PC_reg_N12, ZN 
                           => addr_to_iram_19_port);
   U4394 : TINV_X1 port map( I => n7667, EN => pipeline_stageF_PC_reg_N11, ZN 
                           => addr_to_iram_20_port);
   U4395 : TINV_X1 port map( I => n7668, EN => pipeline_stageF_PC_reg_N10, ZN 
                           => addr_to_iram_21_port);
   U4396 : TINV_X1 port map( I => n7669, EN => pipeline_stageF_PC_reg_N9, ZN =>
                           addr_to_iram_22_port);
   U4397 : TINV_X1 port map( I => n7670, EN => pipeline_stageF_PC_reg_N8, ZN =>
                           addr_to_iram_23_port);
   U4398 : TINV_X1 port map( I => n7671, EN => pipeline_stageF_PC_reg_N7, ZN =>
                           addr_to_iram_24_port);
   U4399 : TINV_X1 port map( I => n7672, EN => pipeline_stageF_PC_reg_N6, ZN =>
                           addr_to_iram_25_port);
   U4400 : TINV_X1 port map( I => n7673, EN => pipeline_stageF_PC_reg_N5, ZN =>
                           addr_to_iram_26_port);
   U4401 : TINV_X1 port map( I => n7674, EN => pipeline_stageF_PC_reg_N4, ZN =>
                           addr_to_iram_27_port);
   U4402 : TINV_X1 port map( I => n7675, EN => pipeline_stageF_PC_reg_N3, ZN =>
                           addr_to_iram_28_port);
   U4403 : TINV_X1 port map( I => n7709, EN => pipeline_stageF_PC_reg_N2, ZN =>
                           addr_to_iram_29_port);
   U4404 : TINV_X1 port map( I => n7710, EN => pipeline_stageF_PC_reg_N1, ZN =>
                           addr_to_iram_30_port);
   pipeline_EXMEM_stage_Forward_sw1_mux_reg : DFF_X1 port map( D => 
                           pipeline_EXMEM_stage_N76, CK => Clk, Q => 
                           pipeline_Forward_sw1_mux, QN => n17380);
   pipeline_MEMWB_Stage_RegDst_Addr_out_MEMWB_reg_4_inst : DFF_X1 port map( D 
                           => pipeline_MEMWB_Stage_N47, CK => Clk, Q => 
                           pipeline_RegDst_to_WB_4_port, QN => n17386);
   pipeline_MEMWB_Stage_RegDst_Addr_out_MEMWB_reg_1_inst : DFF_X1 port map( D 
                           => pipeline_MEMWB_Stage_N44, CK => Clk, Q => 
                           pipeline_RegDst_to_WB_1_port, QN => n17304);
   pipeline_IDEX_Stage_Reg2_Addr_out_IDEX_reg_1_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N204, CK => Clk, Q => 
                           pipeline_Reg2_Addr_to_exe_1_port, QN => net214705);
   pipeline_IDEX_Stage_Reg1_Addr_out_IDEX_reg_0_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N198, CK => Clk, Q => 
                           pipeline_Reg1_Addr_to_exe_0_port, QN => net214704);
   pipeline_IFID_stage_PC_out_IFID_reg_27_inst : DFF_X1 port map( D => n3909, 
                           CK => Clk, Q => pipeline_nextPC_IFID_DEC_27_port, QN
                           => n17469);
   pipeline_IFID_stage_PC_out_IFID_reg_26_inst : DFF_X1 port map( D => n3907, 
                           CK => Clk, Q => pipeline_nextPC_IFID_DEC_26_port, QN
                           => n17466);
   pipeline_IFID_stage_PC_out_IFID_reg_25_inst : DFF_X1 port map( D => n3905, 
                           CK => Clk, Q => pipeline_nextPC_IFID_DEC_25_port, QN
                           => n17451);
   pipeline_IFID_stage_PC_out_IFID_reg_24_inst : DFF_X1 port map( D => n3903, 
                           CK => Clk, Q => pipeline_nextPC_IFID_DEC_24_port, QN
                           => n17465);
   pipeline_IFID_stage_PC_out_IFID_reg_23_inst : DFF_X1 port map( D => n3901, 
                           CK => Clk, Q => pipeline_nextPC_IFID_DEC_23_port, QN
                           => n17435);
   pipeline_IFID_stage_PC_out_IFID_reg_22_inst : DFF_X1 port map( D => n3899, 
                           CK => Clk, Q => pipeline_nextPC_IFID_DEC_22_port, QN
                           => n17464);
   pipeline_IFID_stage_PC_out_IFID_reg_21_inst : DFF_X1 port map( D => n3897, 
                           CK => Clk, Q => pipeline_nextPC_IFID_DEC_21_port, QN
                           => n17448);
   pipeline_IFID_stage_PC_out_IFID_reg_20_inst : DFF_X1 port map( D => n3895, 
                           CK => Clk, Q => pipeline_nextPC_IFID_DEC_20_port, QN
                           => n17463);
   pipeline_IFID_stage_PC_out_IFID_reg_19_inst : DFF_X1 port map( D => n3893, 
                           CK => Clk, Q => pipeline_nextPC_IFID_DEC_19_port, QN
                           => n17438);
   pipeline_IFID_stage_PC_out_IFID_reg_18_inst : DFF_X1 port map( D => n3891, 
                           CK => Clk, Q => pipeline_nextPC_IFID_DEC_18_port, QN
                           => n17462);
   pipeline_IFID_stage_PC_out_IFID_reg_17_inst : DFF_X1 port map( D => n3889, 
                           CK => Clk, Q => pipeline_nextPC_IFID_DEC_17_port, QN
                           => n17443);
   pipeline_IFID_stage_PC_out_IFID_reg_15_inst : DFF_X1 port map( D => n3887, 
                           CK => Clk, Q => pipeline_nextPC_IFID_DEC_15_port, QN
                           => n17453);
   pipeline_IFID_stage_PC_out_IFID_reg_14_inst : DFF_X1 port map( D => n3885, 
                           CK => Clk, Q => pipeline_nextPC_IFID_DEC_14_port, QN
                           => n17460);
   pipeline_IFID_stage_PC_out_IFID_reg_13_inst : DFF_X1 port map( D => n3883, 
                           CK => Clk, Q => pipeline_nextPC_IFID_DEC_13_port, QN
                           => n17442);
   pipeline_IFID_stage_PC_out_IFID_reg_12_inst : DFF_X1 port map( D => n3861, 
                           CK => Clk, Q => pipeline_nextPC_IFID_DEC_12_port, QN
                           => n17459);
   pipeline_IFID_stage_PC_out_IFID_reg_11_inst : DFF_X1 port map( D => n3867, 
                           CK => Clk, Q => pipeline_nextPC_IFID_DEC_11_port, QN
                           => n17441);
   pipeline_IFID_stage_PC_out_IFID_reg_10_inst : DFF_X1 port map( D => n3863, 
                           CK => Clk, Q => pipeline_nextPC_IFID_DEC_10_port, QN
                           => n17458);
   pipeline_IFID_stage_PC_out_IFID_reg_9_inst : DFF_X1 port map( D => n3865, CK
                           => Clk, Q => pipeline_nextPC_IFID_DEC_9_port, QN => 
                           n17436);
   pipeline_IFID_stage_PC_out_IFID_reg_8_inst : DFF_X1 port map( D => n3881, CK
                           => Clk, Q => pipeline_nextPC_IFID_DEC_8_port, QN => 
                           n17457);
   pipeline_IFID_stage_PC_out_IFID_reg_7_inst : DFF_X1 port map( D => n3875, CK
                           => Clk, Q => pipeline_nextPC_IFID_DEC_7_port, QN => 
                           n17468);
   pipeline_IFID_stage_PC_out_IFID_reg_6_inst : DFF_X1 port map( D => n3869, CK
                           => Clk, Q => pipeline_nextPC_IFID_DEC_6_port, QN => 
                           n17456);
   pipeline_IFID_stage_PC_out_IFID_reg_5_inst : DFF_X1 port map( D => n3871, CK
                           => Clk, Q => pipeline_nextPC_IFID_DEC_5_port, QN => 
                           n17454);
   pipeline_IFID_stage_PC_out_IFID_reg_4_inst : DFF_X1 port map( D => n3873, CK
                           => Clk, Q => pipeline_nextPC_IFID_DEC_4_port, QN => 
                           n17455);
   pipeline_IFID_stage_PC_out_IFID_reg_3_inst : DFF_X1 port map( D => n3877, CK
                           => Clk, Q => pipeline_nextPC_IFID_DEC_3_port, QN => 
                           n17439);
   pipeline_IFID_stage_PC_out_IFID_reg_2_inst : DFF_X1 port map( D => n3859, CK
                           => Clk, Q => pipeline_nextPC_IFID_DEC_2_port, QN => 
                           n17470);
   pipeline_IFID_stage_Instr_out_IFID_reg_31_inst : DFF_X1 port map( D => n3957
                           , CK => Clk, Q => pipeline_inst_IFID_DEC_31_port, QN
                           => n17532);
   pipeline_IFID_stage_Instr_out_IFID_reg_23_inst : DFF_X1 port map( D => n3965
                           , CK => Clk, Q => 
                           pipeline_stageD_offset_jump_sign_ext_23_port, QN => 
                           n17383);
   pipeline_EXMEM_stage_ALUres_MEMaddr_out_EXMEM_reg_11_inst : DFF_X1 port map(
                           D => pipeline_EXMEM_stage_N18, CK => Clk, Q => 
                           pipeline_Alu_Out_Addr_to_mem_11_port, QN => 
                           net214703);
   pipeline_EXMEM_stage_ALUres_MEMaddr_out_EXMEM_reg_9_inst : DFF_X1 port map( 
                           D => pipeline_EXMEM_stage_N16, CK => Clk, Q => 
                           pipeline_Alu_Out_Addr_to_mem_9_port, QN => net214702
                           );
   pipeline_EXMEM_stage_ALUres_MEMaddr_out_EXMEM_reg_10_inst : DFF_X1 port map(
                           D => pipeline_EXMEM_stage_N17, CK => Clk, Q => 
                           pipeline_Alu_Out_Addr_to_mem_10_port, QN => 
                           net214701);
   pipeline_EXMEM_stage_ALUres_MEMaddr_out_EXMEM_reg_8_inst : DFF_X1 port map( 
                           D => pipeline_EXMEM_stage_N15, CK => Clk, Q => 
                           pipeline_Alu_Out_Addr_to_mem_8_port, QN => net214700
                           );
   pipeline_EXMEM_stage_ALUres_MEMaddr_out_EXMEM_reg_2_inst : DFF_X1 port map( 
                           D => pipeline_EXMEM_stage_N9, CK => Clk, Q => 
                           pipeline_Alu_Out_Addr_to_mem_2_port, QN => n17398);
   pipeline_IFID_stage_PC_out_IFID_reg_28_inst : DFF_X1 port map( D => n3911, 
                           CK => Clk, Q => pipeline_nextPC_IFID_DEC_28_port, QN
                           => n17467);
   pipeline_EXMEM_stage_ALUres_MEMaddr_out_EXMEM_reg_1_inst : DFF_X1 port map( 
                           D => pipeline_EXMEM_stage_N8, CK => Clk, Q => 
                           pipeline_Alu_Out_Addr_to_mem_1_port, QN => n17397);
   pipeline_EXMEM_stage_ALUres_MEMaddr_out_EXMEM_reg_5_inst : DFF_X1 port map( 
                           D => pipeline_EXMEM_stage_N12, CK => Clk, Q => 
                           pipeline_Alu_Out_Addr_to_mem_5_port, QN => net214699
                           );
   pipeline_EXMEM_stage_ALUres_MEMaddr_out_EXMEM_reg_6_inst : DFF_X1 port map( 
                           D => pipeline_EXMEM_stage_N13, CK => Clk, Q => 
                           pipeline_Alu_Out_Addr_to_mem_6_port, QN => net214698
                           );
   pipeline_EXMEM_stage_ALUres_MEMaddr_out_EXMEM_reg_4_inst : DFF_X1 port map( 
                           D => pipeline_EXMEM_stage_N11, CK => Clk, Q => 
                           pipeline_Alu_Out_Addr_to_mem_4_port, QN => net214697
                           );
   pipeline_EXMEM_stage_ALUres_MEMaddr_out_EXMEM_reg_3_inst : DFF_X1 port map( 
                           D => pipeline_EXMEM_stage_N10, CK => Clk, Q => 
                           pipeline_Alu_Out_Addr_to_mem_3_port, QN => net214696
                           );
   pipeline_EXMEM_stage_ALUres_MEMaddr_out_EXMEM_reg_13_inst : DFF_X1 port map(
                           D => pipeline_EXMEM_stage_N20, CK => Clk, Q => 
                           pipeline_Alu_Out_Addr_to_mem_13_port, QN => 
                           net214695);
   pipeline_IFID_stage_PC_out_IFID_reg_29_inst : DFF_X1 port map( D => n3856, 
                           CK => Clk, Q => pipeline_nextPC_IFID_DEC_29_port, QN
                           => n17452);
   pipeline_EXMEM_stage_ALUres_MEMaddr_out_EXMEM_reg_14_inst : DFF_X1 port map(
                           D => pipeline_EXMEM_stage_N21, CK => Clk, Q => 
                           pipeline_Alu_Out_Addr_to_mem_14_port, QN => 
                           net214694);
   pipeline_IFID_stage_PC_out_IFID_reg_30_inst : DFF_X1 port map( D => n3855, 
                           CK => Clk, Q => pipeline_nextPC_IFID_DEC_30_port, QN
                           => n17471);
   pipeline_EXMEM_stage_ALUres_MEMaddr_out_EXMEM_reg_16_inst : DFF_X1 port map(
                           D => pipeline_EXMEM_stage_N23, CK => Clk, Q => 
                           pipeline_Alu_Out_Addr_to_mem_16_port, QN => 
                           net214693);
   pipeline_EXMEM_stage_ALUres_MEMaddr_out_EXMEM_reg_15_inst : DFF_X1 port map(
                           D => pipeline_EXMEM_stage_N22, CK => Clk, Q => 
                           pipeline_Alu_Out_Addr_to_mem_15_port, QN => 
                           net214692);
   pipeline_EXMEM_stage_ALUres_MEMaddr_out_EXMEM_reg_17_inst : DFF_X1 port map(
                           D => pipeline_EXMEM_stage_N24, CK => Clk, Q => 
                           pipeline_Alu_Out_Addr_to_mem_17_port, QN => 
                           net214691);
   pipeline_EXMEM_stage_ALUres_MEMaddr_out_EXMEM_reg_22_inst : DFF_X1 port map(
                           D => pipeline_EXMEM_stage_N29, CK => Clk, Q => 
                           pipeline_Alu_Out_Addr_to_mem_22_port, QN => 
                           net214690);
   pipeline_EXMEM_stage_ALUres_MEMaddr_out_EXMEM_reg_20_inst : DFF_X1 port map(
                           D => pipeline_EXMEM_stage_N27, CK => Clk, Q => 
                           pipeline_Alu_Out_Addr_to_mem_20_port, QN => 
                           net214689);
   pipeline_EXMEM_stage_ALUres_MEMaddr_out_EXMEM_reg_21_inst : DFF_X1 port map(
                           D => pipeline_EXMEM_stage_N28, CK => Clk, Q => 
                           pipeline_Alu_Out_Addr_to_mem_21_port, QN => 
                           net214688);
   pipeline_EXMEM_stage_ALUres_MEMaddr_out_EXMEM_reg_19_inst : DFF_X1 port map(
                           D => pipeline_EXMEM_stage_N26, CK => Clk, Q => 
                           pipeline_Alu_Out_Addr_to_mem_19_port, QN => 
                           net214687);
   pipeline_EXMEM_stage_ALUres_MEMaddr_out_EXMEM_reg_23_inst : DFF_X1 port map(
                           D => pipeline_EXMEM_stage_N30, CK => Clk, Q => 
                           pipeline_Alu_Out_Addr_to_mem_23_port, QN => 
                           net214686);
   pipeline_EXMEM_stage_ALUres_MEMaddr_out_EXMEM_reg_18_inst : DFF_X1 port map(
                           D => pipeline_EXMEM_stage_N25, CK => Clk, Q => 
                           pipeline_Alu_Out_Addr_to_mem_18_port, QN => 
                           net214685);
   pipeline_EXMEM_stage_ALUres_MEMaddr_out_EXMEM_reg_25_inst : DFF_X1 port map(
                           D => pipeline_EXMEM_stage_N32, CK => Clk, Q => 
                           pipeline_Alu_Out_Addr_to_mem_25_port, QN => 
                           net214684);
   pipeline_EXMEM_stage_ALUres_MEMaddr_out_EXMEM_reg_26_inst : DFF_X1 port map(
                           D => pipeline_EXMEM_stage_N33, CK => Clk, Q => 
                           pipeline_Alu_Out_Addr_to_mem_26_port, QN => 
                           net214683);
   pipeline_EXMEM_stage_ALUres_MEMaddr_out_EXMEM_reg_24_inst : DFF_X1 port map(
                           D => pipeline_EXMEM_stage_N31, CK => Clk, Q => 
                           pipeline_Alu_Out_Addr_to_mem_24_port, QN => 
                           net214682);
   pipeline_EXMEM_stage_ALUres_MEMaddr_out_EXMEM_reg_27_inst : DFF_X1 port map(
                           D => pipeline_EXMEM_stage_N34, CK => Clk, Q => 
                           pipeline_Alu_Out_Addr_to_mem_27_port, QN => 
                           net214681);
   pipeline_EXMEM_stage_ALUres_MEMaddr_out_EXMEM_reg_28_inst : DFF_X1 port map(
                           D => pipeline_EXMEM_stage_N35, CK => Clk, Q => 
                           pipeline_Alu_Out_Addr_to_mem_28_port, QN => 
                           net214680);
   pipeline_EXMEM_stage_ALUres_MEMaddr_out_EXMEM_reg_29_inst : DFF_X1 port map(
                           D => pipeline_EXMEM_stage_N36, CK => Clk, Q => 
                           pipeline_Alu_Out_Addr_to_mem_29_port, QN => 
                           net214679);
   pipeline_EXMEM_stage_ALUres_MEMaddr_out_EXMEM_reg_30_inst : DFF_X1 port map(
                           D => pipeline_EXMEM_stage_N37, CK => Clk, Q => 
                           pipeline_Alu_Out_Addr_to_mem_30_port, QN => 
                           net214678);
   pipeline_EXMEM_stage_ALUres_MEMaddr_out_EXMEM_reg_31_inst : DFF_X1 port map(
                           D => pipeline_EXMEM_stage_N38, CK => Clk, Q => 
                           pipeline_Alu_Out_Addr_to_mem_31_port, QN => 
                           net214677);
   pipeline_IFID_stage_PC_out_IFID_reg_1_inst : DFF_X1 port map( D => n3857, CK
                           => Clk, Q => pipeline_nextPC_IFID_DEC_1_port, QN => 
                           n17446);
   pipeline_IDEX_Stage_Reg2_Addr_out_IDEX_reg_4_inst : DFF_X1 port map( D => 
                           pipeline_IDEX_Stage_N207, CK => Clk, Q => 
                           pipeline_Reg2_Addr_to_exe_4_port, QN => n12625);
   pipeline_EXMEM_stage_RegDst_Addr_out_EXMEM_reg_0_inst : DFF_X1 port map( D 
                           => pipeline_EXMEM_stage_N71, CK => Clk, Q => 
                           pipeline_regDst_to_mem_0_port, QN => n17644);
   pipeline_EXMEM_stage_RegDst_Addr_out_EXMEM_reg_3_inst : DFF_X1 port map( D 
                           => pipeline_EXMEM_stage_N74, CK => Clk, Q => 
                           pipeline_regDst_to_mem_3_port, QN => n17340);
   pipeline_EXMEM_stage_RegDst_Addr_out_EXMEM_reg_4_inst : DFF_X1 port map( D 
                           => pipeline_EXMEM_stage_N75, CK => Clk, Q => 
                           pipeline_regDst_to_mem_4_port, QN => n17393);
   pipeline_EXMEM_stage_ALUres_MEMaddr_out_EXMEM_reg_0_inst : DFF_X1 port map( 
                           D => pipeline_EXMEM_stage_N7, CK => Clk, Q => 
                           pipeline_Alu_Out_Addr_to_mem_0_port, QN => net214676
                           );
   pipeline_IFID_stage_Instr_out_IFID_reg_4_inst : DFF_X1 port map( D => n3983,
                           CK => Clk, Q => 
                           pipeline_stageD_offset_to_jump_temp_4_port, QN => 
                           n17412);
   U11979 : NAND3_X1 port map( A1 => n13980, A2 => n17704, A3 => n13984, ZN => 
                           pipeline_cu_pipeline_N107);
   U11980 : NAND3_X1 port map( A1 => n14028, A2 => n14019, A3 => n14029, ZN => 
                           n14027);
   U11981 : NAND3_X1 port map( A1 => pipeline_inst_IFID_DEC_29_port, A2 => 
                           n13995, A3 => n17348, ZN => n14035);
   U11982 : NAND3_X1 port map( A1 => n14005, A2 => n14044, A3 => n14032, ZN => 
                           n14021);
   U11983 : NAND3_X1 port map( A1 => n14049, A2 => n14000, A3 => n17382, ZN => 
                           n14048);
   U11984 : NAND3_X1 port map( A1 => n14000, A2 => n17348, A3 => 
                           pipeline_inst_IFID_DEC_29_port, ZN => n14070);
   U11985 : NAND3_X1 port map( A1 => pipeline_WB_controls_in_MEMWB_1_port, A2 
                           => pipeline_MEM_controls_in_MEM_1_port, A3 => n14090
                           , ZN => n14089);
   U11986 : NAND3_X1 port map( A1 => pipeline_WB_controls_in_EXMEM_1_port, A2 
                           => pipeline_MEM_controls_in_EXMEM_1_port, A3 => 
                           n14095, ZN => n14086);
   U11987 : XOR2_X1 port map( A => n17384, B => n14100, Z => n14099);
   U11988 : XOR2_X1 port map( A => n17328, B => n14101, Z => n14097);
   U11993 : XOR2_X1 port map( A => n17383, B => n14113, Z => n14098);
   U11994 : NAND3_X1 port map( A1 => pipeline_WB_controls_in_EXMEM_1_port, A2 
                           => pipeline_MEM_controls_in_EXMEM_1_port, A3 => 
                           n13983, ZN => n14094);
   U11995 : NAND3_X1 port map( A1 => pipeline_cu_pipeline_N89, A2 => n17428, A3
                           => n17361, ZN => n14174);
   U11996 : NAND3_X1 port map( A1 => pipeline_stageD_offset_to_jump_temp_5_port
                           , A2 => n14067, A3 => n17406, ZN => n14066);
   U11997 : NAND3_X1 port map( A1 => pipeline_inst_IFID_DEC_29_port, A2 => 
                           n14049, A3 => n17313, ZN => n14058);
   U11998 : NAND3_X1 port map( A1 => pipeline_inst_IFID_DEC_27_port, A2 => 
                           n14001, A3 => n17347, ZN => n14029);
   U11999 : NAND3_X1 port map( A1 => pipeline_inst_IFID_DEC_31_port, A2 => 
                           n14084, A3 => n17348, ZN => n14169);
   U12000 : NAND3_X1 port map( A1 => n14241, A2 => n14242, A3 => n14243, ZN => 
                           n14201);
   U12001 : NAND3_X1 port map( A1 => n14268, A2 => n14269, A3 => n14270, ZN => 
                           n14252);
   U12002 : NAND3_X1 port map( A1 => n14288, A2 => n14289, A3 => n14290, ZN => 
                           n14272);
   U12003 : NAND3_X1 port map( A1 => n14308, A2 => n14309, A3 => n14310, ZN => 
                           n14292);
   U12004 : NAND3_X1 port map( A1 => n14328, A2 => n14329, A3 => n14330, ZN => 
                           n14312);
   U12005 : NAND3_X1 port map( A1 => n14348, A2 => n14349, A3 => n14350, ZN => 
                           n14332);
   U12006 : NAND3_X1 port map( A1 => n14368, A2 => n14369, A3 => n14370, ZN => 
                           n14352);
   U12007 : NAND3_X1 port map( A1 => n14388, A2 => n14389, A3 => n14390, ZN => 
                           n14372);
   U12008 : NAND3_X1 port map( A1 => n14408, A2 => n14409, A3 => n14410, ZN => 
                           n14392);
   U12009 : NAND3_X1 port map( A1 => n14428, A2 => n14429, A3 => n14430, ZN => 
                           n14412);
   U12010 : NAND3_X1 port map( A1 => n14448, A2 => n14449, A3 => n14450, ZN => 
                           n14432);
   U12011 : NAND3_X1 port map( A1 => n14468, A2 => n14469, A3 => n14470, ZN => 
                           n14452);
   U12012 : NAND3_X1 port map( A1 => n14488, A2 => n14489, A3 => n14490, ZN => 
                           n14472);
   U12013 : NAND3_X1 port map( A1 => n14508, A2 => n14509, A3 => n14510, ZN => 
                           n14492);
   U12014 : NAND3_X1 port map( A1 => n14528, A2 => n14529, A3 => n14530, ZN => 
                           n14512);
   U12015 : NAND3_X1 port map( A1 => n14548, A2 => n14549, A3 => n14550, ZN => 
                           n14532);
   U12016 : NAND3_X1 port map( A1 => n14568, A2 => n14569, A3 => n14570, ZN => 
                           n14552);
   U12017 : NAND3_X1 port map( A1 => n14588, A2 => n14589, A3 => n14590, ZN => 
                           n14572);
   U12018 : NAND3_X1 port map( A1 => n14608, A2 => n14609, A3 => n14610, ZN => 
                           n14592);
   U12019 : NAND3_X1 port map( A1 => n14628, A2 => n14629, A3 => n14630, ZN => 
                           n14612);
   U12020 : NAND3_X1 port map( A1 => n14648, A2 => n14649, A3 => n14650, ZN => 
                           n14632);
   U12021 : NAND3_X1 port map( A1 => n14668, A2 => n14669, A3 => n14670, ZN => 
                           n14652);
   U12022 : NAND3_X1 port map( A1 => n14688, A2 => n14689, A3 => n14690, ZN => 
                           n14672);
   U12023 : NAND3_X1 port map( A1 => n14708, A2 => n14709, A3 => n14710, ZN => 
                           n14692);
   U12024 : NAND3_X1 port map( A1 => n14728, A2 => n14729, A3 => n14730, ZN => 
                           n14712);
   U12025 : NAND3_X1 port map( A1 => n14748, A2 => n14749, A3 => n14750, ZN => 
                           n14732);
   U12026 : NAND3_X1 port map( A1 => n14768, A2 => n14769, A3 => n14770, ZN => 
                           n14752);
   U12027 : NAND3_X1 port map( A1 => n14788, A2 => n14789, A3 => n14790, ZN => 
                           n14772);
   U12028 : NAND3_X1 port map( A1 => n14808, A2 => n14809, A3 => n14810, ZN => 
                           n14792);
   U12029 : NAND3_X1 port map( A1 => n14828, A2 => n14829, A3 => n14830, ZN => 
                           n14812);
   U12030 : NAND3_X1 port map( A1 => n14848, A2 => n14849, A3 => n14850, ZN => 
                           n14832);
   U12031 : NAND3_X1 port map( A1 => 
                           pipeline_stageD_offset_jump_sign_ext_16_port, A2 => 
                           n17407, A3 => n17349, ZN => n14861);
   U12032 : NAND3_X1 port map( A1 => 
                           pipeline_stageD_offset_jump_sign_ext_19_port, A2 => 
                           pipeline_stageD_offset_jump_sign_ext_16_port, A3 => 
                           n17407, ZN => n14867);
   U12033 : NAND3_X1 port map( A1 => 
                           pipeline_stageD_offset_jump_sign_ext_19_port, A2 => 
                           n17407, A3 => n17316, ZN => n14866);
   U12034 : NAND3_X1 port map( A1 => 
                           pipeline_stageD_offset_jump_sign_ext_20_port, A2 => 
                           n17349, A3 => n17316, ZN => n14872);
   U12035 : NAND3_X1 port map( A1 => 
                           pipeline_stageD_offset_jump_sign_ext_20_port, A2 => 
                           pipeline_stageD_offset_jump_sign_ext_16_port, A3 => 
                           n17349, ZN => n14873);
   U12036 : NAND3_X1 port map( A1 => n14880, A2 => n14881, A3 => n14882, ZN => 
                           n14852);
   U12037 : NAND3_X1 port map( A1 => n17407, A2 => n17349, A3 => n17316, ZN => 
                           n14862);
   U12038 : NAND3_X1 port map( A1 => 
                           pipeline_stageD_offset_jump_sign_ext_19_port, A2 => 
                           pipeline_stageD_offset_jump_sign_ext_20_port, A3 => 
                           n17316, ZN => n14878);
   U12039 : NAND3_X1 port map( A1 => 
                           pipeline_stageD_offset_jump_sign_ext_20_port, A2 => 
                           pipeline_stageD_offset_jump_sign_ext_19_port, A3 => 
                           pipeline_stageD_offset_jump_sign_ext_16_port, ZN => 
                           n14879);
   U12040 : NAND3_X1 port map( A1 => n14952, A2 => n12649, A3 => n17740, ZN => 
                           n14951);
   U12041 : NAND3_X1 port map( A1 => n14958, A2 => n14959, A3 => n14960, ZN => 
                           n14957);
   U12042 : OAI33_X1 port map( A1 => n17074, A2 => n14967, A3 => n12649, B1 => 
                           n17740, B2 => n14968, B3 => n17091, ZN => n14956);
   U12043 : NAND3_X1 port map( A1 => n17103, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_1_port, A3 
                           => n14954, ZN => n14972);
   U12044 : NAND3_X1 port map( A1 => n14977, A2 => n14978, A3 => n14979, ZN => 
                           n14976);
   U12045 : MUX2_X1 port map( A => n13934, B => n13929, S => n17430, Z => 
                           n14120);
   U12046 : NAND3_X1 port map( A1 => n17104, A2 => n15133, A3 => n14954, ZN => 
                           n15131);
   U12047 : OAI33_X1 port map( A1 => n15133, A2 => n17679, A3 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N136, B1 => n15134
                           , B2 => n14968, B3 => n17104, ZN => n15126);
   U12050 : NAND3_X1 port map( A1 => pipeline_stageE_EXE_ALU_alu_shift_N136, A2
                           => n14952, A3 => n15134, ZN => n15124);
   U12051 : NAND3_X1 port map( A1 => n14952, A2 => 
                           pipeline_stageE_input1_to_ALU_30_port, A3 => n15150,
                           ZN => n15149);
   U12052 : NAND3_X1 port map( A1 => n15154, A2 => n15155, A3 => n15156, ZN => 
                           n15153);
   U12053 : OAI33_X1 port map( A1 => n15157, A2 => n17678, A3 => 
                           pipeline_stageE_input1_to_ALU_30_port, B1 => n15150,
                           B2 => n14968, B3 => n17083, ZN => n15152);
   U12054 : XOR2_X1 port map( A => n15159, B => n15160, Z => n15009);
   U12055 : NAND3_X1 port map( A1 => n14952, A2 => 
                           pipeline_stageE_input1_to_ALU_29_port, A3 => n15169,
                           ZN => n15168);
   U12056 : NAND3_X1 port map( A1 => n15173, A2 => n15174, A3 => n15175, ZN => 
                           n15172);
   U12057 : OAI33_X1 port map( A1 => n15176, A2 => n14967, A3 => 
                           pipeline_stageE_input1_to_ALU_29_port, B1 => n15169,
                           B2 => n14968, B3 => n17094, ZN => n15171);
   U12058 : NAND3_X1 port map( A1 => n14952, A2 => 
                           pipeline_stageE_input1_to_ALU_28_port, A3 => n15182,
                           ZN => n15181);
   U12059 : NAND3_X1 port map( A1 => n15186, A2 => n15187, A3 => n15188, ZN => 
                           n15185);
   U12060 : OAI33_X1 port map( A1 => n15189, A2 => n17679, A3 => 
                           pipeline_stageE_input1_to_ALU_28_port, B1 => n15182,
                           B2 => n14968, B3 => n17093, ZN => n15184);
   U12061 : NAND3_X1 port map( A1 => n17078, A2 => n15201, A3 => n14954, ZN => 
                           n15199);
   U12062 : OAI33_X1 port map( A1 => n15201, A2 => n17678, A3 => 
                           pipeline_stageE_input1_to_ALU_27_port, B1 => n15202,
                           B2 => n14968, B3 => n17078, ZN => n15194);
   U12064 : NAND3_X1 port map( A1 => pipeline_stageE_input1_to_ALU_27_port, A2 
                           => n14952, A3 => n15202, ZN => n15192);
   U12065 : NAND3_X1 port map( A1 => n17086, A2 => n15215, A3 => n14954, ZN => 
                           n15213);
   U12066 : OAI33_X1 port map( A1 => n15215, A2 => n14967, A3 => 
                           pipeline_stageE_input1_to_ALU_26_port, B1 => n15216,
                           B2 => n14968, B3 => n17086, ZN => n15208);
   U12067 : NAND3_X1 port map( A1 => pipeline_stageE_input1_to_ALU_26_port, A2 
                           => n14952, A3 => n15216, ZN => n15206);
   U12068 : NAND3_X1 port map( A1 => n14952, A2 => n17159, A3 => n15224, ZN => 
                           n15223);
   U12069 : NAND3_X1 port map( A1 => n15228, A2 => n15229, A3 => n15230, ZN => 
                           n15227);
   U12070 : OAI33_X1 port map( A1 => n15231, A2 => n17679, A3 => n17159, B1 => 
                           n15224, B2 => n14968, B3 => n17115, ZN => n15226);
   U12071 : NAND3_X1 port map( A1 => n17117, A2 => n15245, A3 => n14954, ZN => 
                           n15243);
   U12072 : OAI33_X1 port map( A1 => n15245, A2 => n17678, A3 => n17158, B1 => 
                           n15246, B2 => n14968, B3 => n17117, ZN => n15238);
   U12073 : XOR2_X1 port map( A => n15247, B => n15248, Z => n15013);
   U12074 : NAND3_X1 port map( A1 => n17158, A2 => n14952, A3 => n15246, ZN => 
                           n15236);
   U12075 : NAND3_X1 port map( A1 => n17092, A2 => n15260, A3 => n17677, ZN => 
                           n15258);
   U12076 : OAI33_X1 port map( A1 => n15260, A2 => n14967, A3 => 
                           pipeline_stageE_input1_to_ALU_23_port, B1 => n15261,
                           B2 => n14968, B3 => n17092, ZN => n15253);
   U12077 : XOR2_X1 port map( A => n15262, B => n15263, Z => n15022);
   U12078 : NAND3_X1 port map( A1 => pipeline_stageE_input1_to_ALU_23_port, A2 
                           => n14952, A3 => n15261, ZN => n15251);
   U12079 : NAND3_X1 port map( A1 => n17116, A2 => n15278, A3 => n17677, ZN => 
                           n15276);
   U12080 : OAI33_X1 port map( A1 => n15278, A2 => n17679, A3 => 
                           pipeline_stageE_input1_to_ALU_22_port, B1 => n15279,
                           B2 => n14968, B3 => n17116, ZN => n15271);
   U12081 : NAND3_X1 port map( A1 => pipeline_stageE_input1_to_ALU_22_port, A2 
                           => n14952, A3 => n15279, ZN => n15269);
   U12082 : NAND3_X1 port map( A1 => n14952, A2 => 
                           pipeline_stageE_input1_to_ALU_21_port, A3 => n15285,
                           ZN => n15284);
   U12083 : NAND3_X1 port map( A1 => n15289, A2 => n15290, A3 => n15291, ZN => 
                           n15288);
   U12084 : OAI33_X1 port map( A1 => n15292, A2 => n17678, A3 => 
                           pipeline_stageE_input1_to_ALU_21_port, B1 => n15285,
                           B2 => n14968, B3 => n17084, ZN => n15287);
   U12085 : XOR2_X1 port map( A => n15294, B => n15295, Z => n15017);
   U12086 : NAND3_X1 port map( A1 => n17118, A2 => n15311, A3 => n17677, ZN => 
                           n15309);
   U12087 : OAI33_X1 port map( A1 => n15311, A2 => n14967, A3 => n17157, B1 => 
                           n15312, B2 => n14968, B3 => n17118, ZN => n15304);
   U12088 : NAND3_X1 port map( A1 => n17157, A2 => n14952, A3 => n15312, ZN => 
                           n15302);
   U12089 : NAND3_X1 port map( A1 => n17097, A2 => n15330, A3 => n17677, ZN => 
                           n15328);
   U12090 : OAI33_X1 port map( A1 => n15330, A2 => n17679, A3 => 
                           pipeline_stageE_input1_to_ALU_19_port, B1 => n15331,
                           B2 => n14968, B3 => n17097, ZN => n15323);
   U12091 : XOR2_X1 port map( A => n15332, B => n15333, Z => n15023);
   U12092 : XOR2_X1 port map( A => n15334, B => n17097, Z => n15333);
   U12093 : NAND3_X1 port map( A1 => pipeline_stageE_input1_to_ALU_19_port, A2 
                           => n14952, A3 => n15331, ZN => n15321);
   U12094 : NAND3_X1 port map( A1 => n17096, A2 => n15345, A3 => n17677, ZN => 
                           n15343);
   U12095 : OAI33_X1 port map( A1 => n15345, A2 => n17678, A3 => 
                           pipeline_stageE_input1_to_ALU_18_port, B1 => n15346,
                           B2 => n14968, B3 => n17096, ZN => n15338);
   U12097 : NAND3_X1 port map( A1 => pipeline_stageE_input1_to_ALU_18_port, A2 
                           => n14952, A3 => n15346, ZN => n15336);
   U12098 : NAND3_X1 port map( A1 => n17079, A2 => n15362, A3 => n17677, ZN => 
                           n15360);
   U12099 : OAI33_X1 port map( A1 => n15362, A2 => n14967, A3 => 
                           pipeline_stageE_input1_to_ALU_17_port, B1 => n15363,
                           B2 => n14968, B3 => n17079, ZN => n15355);
   U12101 : NAND3_X1 port map( A1 => pipeline_stageE_input1_to_ALU_17_port, A2 
                           => n14952, A3 => n15363, ZN => n15353);
   U12102 : NAND3_X1 port map( A1 => n14952, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_A_16_port, A3 
                           => n15372, ZN => n15371);
   U12103 : NAND3_X1 port map( A1 => n15376, A2 => n15377, A3 => n15378, ZN => 
                           n15375);
   U12104 : OAI33_X1 port map( A1 => n15379, A2 => n17679, A3 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_A_16_port, B1 
                           => n15372, B2 => n14968, B3 => n17738, ZN => n15374)
                           ;
   U12105 : XOR2_X1 port map( A => n15381, B => n15368, Z => n15032);
   U12106 : NAND3_X1 port map( A1 => n14952, A2 => 
                           pipeline_stageE_input1_to_ALU_15_port, A3 => n15386,
                           ZN => n15385);
   U12107 : NAND3_X1 port map( A1 => n15390, A2 => n15391, A3 => n15392, ZN => 
                           n15389);
   U12108 : OAI33_X1 port map( A1 => n15393, A2 => n17678, A3 => 
                           pipeline_stageE_input1_to_ALU_15_port, B1 => n15386,
                           B2 => n14968, B3 => n17101, ZN => n15388);
   U12109 : XOR2_X1 port map( A => n15395, B => n15396, Z => n15029);
   U12110 : XOR2_X1 port map( A => n17101, B => n15397, Z => n15396);
   U12111 : NAND3_X1 port map( A1 => n17100, A2 => n15410, A3 => n17677, ZN => 
                           n15408);
   U12112 : OAI33_X1 port map( A1 => n15410, A2 => n14967, A3 => 
                           pipeline_stageE_input1_to_ALU_14_port, B1 => n15411,
                           B2 => n14968, B3 => n17100, ZN => n15403);
   U12113 : XOR2_X1 port map( A => n15399, B => n15412, Z => n15027);
   U12114 : NAND3_X1 port map( A1 => pipeline_stageE_input1_to_ALU_14_port, A2 
                           => n14952, A3 => n15411, ZN => n15401);
   U12115 : NAND3_X1 port map( A1 => n15425, A2 => n15426, A3 => n17677, ZN => 
                           n15424);
   U12116 : OAI33_X1 port map( A1 => n15426, A2 => n17679, A3 => n17160, B1 => 
                           n15427, B2 => n14968, B3 => n15425, ZN => n15419);
   U12117 : XOR2_X1 port map( A => n15428, B => n15415, Z => n15033);
   U12118 : NAND3_X1 port map( A1 => n17160, A2 => n14952, A3 => n15427, ZN => 
                           n15417);
   U12119 : NAND3_X1 port map( A1 => n14952, A2 => 
                           pipeline_stageE_input1_to_ALU_12_port, A3 => n15435,
                           ZN => n15434);
   U12120 : NAND3_X1 port map( A1 => n15439, A2 => n15440, A3 => n15441, ZN => 
                           n15438);
   U12121 : OAI33_X1 port map( A1 => n15442, A2 => n17678, A3 => 
                           pipeline_stageE_input1_to_ALU_12_port, B1 => n15435,
                           B2 => n14968, B3 => n17080, ZN => n15437);
   U12122 : XOR2_X1 port map( A => n15444, B => n15429, Z => n15030);
   U12123 : NAND3_X1 port map( A1 => n14952, A2 => 
                           pipeline_stageE_input1_to_ALU_11_port, A3 => n15449,
                           ZN => n15448);
   U12124 : NAND3_X1 port map( A1 => n15453, A2 => n15454, A3 => n15455, ZN => 
                           n15452);
   U12125 : OAI33_X1 port map( A1 => n15456, A2 => n14967, A3 => 
                           pipeline_stageE_input1_to_ALU_11_port, B1 => n15449,
                           B2 => n14968, B3 => n17082, ZN => n15451);
   U12126 : NAND3_X1 port map( A1 => n17085, A2 => n15473, A3 => n14954, ZN => 
                           n15471);
   U12127 : OAI33_X1 port map( A1 => n15473, A2 => n17679, A3 => 
                           pipeline_stageE_input1_to_ALU_10_port, B1 => n15474,
                           B2 => n14968, B3 => n17085, ZN => n15466);
   U12128 : XOR2_X1 port map( A => n15475, B => n15462, Z => n15034);
   U12129 : NAND3_X1 port map( A1 => pipeline_stageE_input1_to_ALU_10_port, A2 
                           => n14952, A3 => n15474, ZN => n15464);
   U12130 : NAND3_X1 port map( A1 => n17090, A2 => n15491, A3 => n14954, ZN => 
                           n15489);
   U12131 : OAI33_X1 port map( A1 => n15491, A2 => n17678, A3 => 
                           pipeline_stageE_input1_to_ALU_9_port, B1 => n15492, 
                           B2 => n14968, B3 => n17090, ZN => n15484);
   U12132 : NAND3_X1 port map( A1 => pipeline_stageE_input1_to_ALU_9_port, A2 
                           => n14952, A3 => n15492, ZN => n15482);
   U12133 : NAND3_X1 port map( A1 => n14952, A2 => 
                           pipeline_stageE_input1_to_ALU_8_port, A3 => n15498, 
                           ZN => n15497);
   U12134 : NAND3_X1 port map( A1 => n15502, A2 => n15503, A3 => n15504, ZN => 
                           n15501);
   U12135 : OAI33_X1 port map( A1 => n15505, A2 => n14967, A3 => 
                           pipeline_stageE_input1_to_ALU_8_port, B1 => n15498, 
                           B2 => n14968, B3 => n17095, ZN => n15500);
   U12136 : XOR2_X1 port map( A => n15507, B => n15508, Z => n15039);
   U12137 : NAND3_X1 port map( A1 => n14952, A2 => 
                           pipeline_stageE_input1_to_ALU_7_port, A3 => n15512, 
                           ZN => n15511);
   U12138 : NAND3_X1 port map( A1 => n15516, A2 => n15517, A3 => n15518, ZN => 
                           n15515);
   U12139 : OAI33_X1 port map( A1 => n15519, A2 => n17679, A3 => 
                           pipeline_stageE_input1_to_ALU_7_port, B1 => n15512, 
                           B2 => n14968, B3 => n17089, ZN => n15514);
   U12140 : NAND3_X1 port map( A1 => n17088, A2 => n15537, A3 => n14954, ZN => 
                           n15535);
   U12141 : OAI33_X1 port map( A1 => n15537, A2 => n17678, A3 => 
                           pipeline_stageE_input1_to_ALU_6_port, B1 => n15538, 
                           B2 => n14968, B3 => n17088, ZN => n15530);
   U12142 : NAND3_X1 port map( A1 => pipeline_stageE_input1_to_ALU_6_port, A2 
                           => n14952, A3 => n15538, ZN => n15528);
   U12143 : NAND3_X1 port map( A1 => n17087, A2 => n15552, A3 => n14954, ZN => 
                           n15550);
   U12144 : OAI33_X1 port map( A1 => n15552, A2 => n14967, A3 => 
                           pipeline_stageE_input1_to_ALU_5_port, B1 => n15553, 
                           B2 => n14968, B3 => n17087, ZN => n15545);
   U12145 : NAND3_X1 port map( A1 => pipeline_stageE_input1_to_ALU_5_port, A2 
                           => n14952, A3 => n15553, ZN => n15543);
   U12146 : NAND3_X1 port map( A1 => n15564, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, A3 
                           => n14954, ZN => n15563);
   U12147 : OAI33_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, A2 
                           => n17679, A3 => 
                           pipeline_stageE_input1_to_ALU_4_port, B1 => n17737, 
                           B2 => n14968, B3 => n15564, ZN => n15558);
   U12148 : XOR2_X1 port map( A => n15566, B => n15567, Z => n15041);
   U12149 : NAND3_X1 port map( A1 => n14952, A2 => n17739, A3 => 
                           pipeline_stageE_input1_to_ALU_3_port, ZN => n15571);
   U12150 : NAND3_X1 port map( A1 => n15577, A2 => n15578, A3 => n15579, ZN => 
                           n15576);
   U12151 : NAND3_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_5_port, 
                           A2 => pipeline_EXE_controls_in_EXEcute_6_port, A3 =>
                           n17705, ZN => n15586);
   U12152 : OAI33_X1 port map( A1 => n17077, A2 => n14968, A3 => n17739, B1 => 
                           pipeline_stageE_input1_to_ALU_3_port, B2 => n17678, 
                           B3 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_3_port, ZN 
                           => n15575);
   U12154 : XOR2_X1 port map( A => n15590, B => n15591, Z => n15045);
   U12155 : MUX2_X1 port map( A => n15592, B => n15593, S => n17381, Z => 
                           n15591);
   U12156 : NAND3_X1 port map( A1 => n15596, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N202, A3 => n15050
                           , ZN => n15595);
   U12157 : XOR2_X1 port map( A => n15598, B => n17077, Z => n15590);
   U12158 : NAND3_X1 port map( A1 => n15602, A2 => n15603, A3 => n15604, ZN => 
                           n3991);
   U12161 : NAND3_X1 port map( A1 => n15689, A2 => n15690, A3 => n15691, ZN => 
                           n3912);
   U12162 : NAND3_X1 port map( A1 => n15694, A2 => n15695, A3 => n15696, ZN => 
                           n3910);
   U12163 : NAND3_X1 port map( A1 => n15699, A2 => n15700, A3 => n15701, ZN => 
                           n3908);
   U12164 : NAND3_X1 port map( A1 => n15704, A2 => n15705, A3 => n15706, ZN => 
                           n3906);
   U12165 : NAND3_X1 port map( A1 => n15709, A2 => n15710, A3 => n15711, ZN => 
                           n3904);
   U12166 : NAND3_X1 port map( A1 => n15714, A2 => n15715, A3 => n15716, ZN => 
                           n3902);
   U12167 : NAND3_X1 port map( A1 => n15719, A2 => n15720, A3 => n15721, ZN => 
                           n3900);
   U12168 : NAND3_X1 port map( A1 => n15724, A2 => n15725, A3 => n15726, ZN => 
                           n3898);
   U12169 : NAND3_X1 port map( A1 => n15729, A2 => n15730, A3 => n15731, ZN => 
                           n3896);
   U12170 : NAND3_X1 port map( A1 => n15734, A2 => n15735, A3 => n15736, ZN => 
                           n3894);
   U12171 : NAND3_X1 port map( A1 => n15739, A2 => n15740, A3 => n15741, ZN => 
                           n3892);
   U12172 : NAND3_X1 port map( A1 => n15744, A2 => n15745, A3 => n15746, ZN => 
                           n3890);
   U12173 : NAND3_X1 port map( A1 => n15749, A2 => n15750, A3 => n15751, ZN => 
                           n3888);
   U12174 : NAND3_X1 port map( A1 => n15754, A2 => n15755, A3 => n15756, ZN => 
                           n3886);
   U12175 : NAND3_X1 port map( A1 => n15759, A2 => n15760, A3 => n15761, ZN => 
                           n3884);
   U12176 : NAND3_X1 port map( A1 => n15764, A2 => n15765, A3 => n15766, ZN => 
                           n3882);
   U12177 : NAND3_X1 port map( A1 => n15769, A2 => n15770, A3 => n15771, ZN => 
                           n3880);
   U12178 : NAND3_X1 port map( A1 => n15774, A2 => n15775, A3 => n15776, ZN => 
                           n3878);
   U12179 : NAND3_X1 port map( A1 => n15779, A2 => n15780, A3 => n15781, ZN => 
                           n3876);
   U12180 : NAND3_X1 port map( A1 => n15784, A2 => n15785, A3 => n15786, ZN => 
                           n3874);
   U12181 : NAND3_X1 port map( A1 => n15789, A2 => n15790, A3 => n15791, ZN => 
                           n3872);
   U12182 : NAND3_X1 port map( A1 => n15794, A2 => n15795, A3 => n15796, ZN => 
                           n3870);
   U12183 : NAND3_X1 port map( A1 => n15799, A2 => n15800, A3 => n15801, ZN => 
                           n3868);
   U12184 : NAND3_X1 port map( A1 => n15804, A2 => n15805, A3 => n15806, ZN => 
                           n3866);
   U12185 : NAND3_X1 port map( A1 => n15809, A2 => n15810, A3 => n15811, ZN => 
                           n3864);
   U12186 : NAND3_X1 port map( A1 => n15814, A2 => n15815, A3 => n15816, ZN => 
                           n3862);
   U12187 : NAND3_X1 port map( A1 => n15819, A2 => n15820, A3 => n15821, ZN => 
                           n3860);
   U12188 : NAND3_X1 port map( A1 => n15824, A2 => n15825, A3 => n15826, ZN => 
                           n3858);
   U12189 : NAND3_X1 port map( A1 => n15839, A2 => n14125, A3 => n15646, ZN => 
                           n15841);
   U12190 : NAND3_X1 port map( A1 => n14049, A2 => n17382, A3 => n17313, ZN => 
                           n14186);
   U12191 : NAND3_X1 port map( A1 => n15844, A2 => n15845, A3 => n15830, ZN => 
                           n15843);
   U12192 : OAI33_X1 port map( A1 => n15887, A2 => n15827, A3 => n15888, B1 => 
                           n15889, B2 => n15890, B3 => n15891, ZN => n15886);
   U12193 : NAND3_X1 port map( A1 => n15932, A2 => n15933, A3 => n15934, ZN => 
                           n15892);
   U12194 : NAND3_X1 port map( A1 => n15958, A2 => n15959, A3 => n15960, ZN => 
                           n15942);
   U12195 : NAND3_X1 port map( A1 => n15977, A2 => n15978, A3 => n15979, ZN => 
                           n15961);
   U12196 : NAND3_X1 port map( A1 => n15996, A2 => n15997, A3 => n15998, ZN => 
                           n15980);
   U12197 : NAND3_X1 port map( A1 => n16021, A2 => n16022, A3 => n16023, ZN => 
                           n16005);
   U12198 : NAND3_X1 port map( A1 => n16040, A2 => n16041, A3 => n16042, ZN => 
                           n16024);
   U12199 : NAND3_X1 port map( A1 => n16059, A2 => n16060, A3 => n16061, ZN => 
                           n16043);
   U12200 : NAND3_X1 port map( A1 => n16078, A2 => n16079, A3 => n16080, ZN => 
                           n16062);
   U12201 : NAND3_X1 port map( A1 => n16097, A2 => n16098, A3 => n16099, ZN => 
                           n16081);
   U12202 : NAND3_X1 port map( A1 => n16116, A2 => n16117, A3 => n16118, ZN => 
                           n16100);
   U12203 : NAND3_X1 port map( A1 => n16135, A2 => n16136, A3 => n16137, ZN => 
                           n16119);
   U12204 : NAND3_X1 port map( A1 => n16154, A2 => n16155, A3 => n16156, ZN => 
                           n16138);
   U12205 : NAND3_X1 port map( A1 => n16173, A2 => n16174, A3 => n16175, ZN => 
                           n16157);
   U12206 : NAND3_X1 port map( A1 => n16192, A2 => n16193, A3 => n16194, ZN => 
                           n16176);
   U12207 : NAND3_X1 port map( A1 => n16211, A2 => n16212, A3 => n16213, ZN => 
                           n16195);
   U12208 : NAND3_X1 port map( A1 => n16230, A2 => n16231, A3 => n16232, ZN => 
                           n16214);
   U12209 : NAND3_X1 port map( A1 => n16249, A2 => n16250, A3 => n16251, ZN => 
                           n16233);
   U12210 : NAND3_X1 port map( A1 => n16268, A2 => n16269, A3 => n16270, ZN => 
                           n16252);
   U12211 : NAND3_X1 port map( A1 => n16287, A2 => n16288, A3 => n16289, ZN => 
                           n16271);
   U12212 : NAND3_X1 port map( A1 => n16306, A2 => n16307, A3 => n16308, ZN => 
                           n16290);
   U12213 : NAND3_X1 port map( A1 => n16326, A2 => n16327, A3 => n16328, ZN => 
                           n16310);
   U12214 : NAND3_X1 port map( A1 => n16345, A2 => n16346, A3 => n16347, ZN => 
                           n16329);
   U12215 : NAND3_X1 port map( A1 => n16364, A2 => n16365, A3 => n16366, ZN => 
                           n16348);
   U12216 : NAND3_X1 port map( A1 => n16383, A2 => n16384, A3 => n16385, ZN => 
                           n16367);
   U12217 : NAND3_X1 port map( A1 => n16398, A2 => n16399, A3 => n16400, ZN => 
                           n16387);
   U12218 : NAND3_X1 port map( A1 => n16417, A2 => n16418, A3 => n16419, ZN => 
                           n16406);
   U12219 : NAND3_X1 port map( A1 => n16440, A2 => n16441, A3 => n16442, ZN => 
                           n16424);
   U12220 : NAND3_X1 port map( A1 => n16459, A2 => n16460, A3 => n16461, ZN => 
                           n16443);
   U12221 : NAND3_X1 port map( A1 => n16478, A2 => n16479, A3 => n16480, ZN => 
                           n16462);
   U12222 : NAND3_X1 port map( A1 => n16497, A2 => n16498, A3 => n16499, ZN => 
                           n16481);
   U12223 : NAND3_X1 port map( A1 => n16516, A2 => n16517, A3 => n16518, ZN => 
                           n16500);
   U12224 : NAND3_X1 port map( A1 => 
                           pipeline_stageD_offset_jump_sign_ext_21_port, A2 => 
                           n17384, A3 => n17328, ZN => n16528);
   U12225 : NAND3_X1 port map( A1 => n17384, A2 => n17328, A3 => n17315, ZN => 
                           n16531);
   U12226 : NAND3_X1 port map( A1 => 
                           pipeline_stageD_offset_jump_sign_ext_24_port, A2 => 
                           pipeline_stageD_offset_jump_sign_ext_21_port, A3 => 
                           n17328, ZN => n16534);
   U12227 : NAND3_X1 port map( A1 => 
                           pipeline_stageD_offset_jump_sign_ext_31_port, A2 => 
                           n17384, A3 => n17315, ZN => n16539);
   U12228 : NAND3_X1 port map( A1 => 
                           pipeline_stageD_offset_jump_sign_ext_31_port, A2 => 
                           pipeline_stageD_offset_jump_sign_ext_21_port, A3 => 
                           n17384, ZN => n16540);
   U12229 : NAND3_X1 port map( A1 => n16547, A2 => n16548, A3 => n16549, ZN => 
                           n16519);
   U12230 : NAND3_X1 port map( A1 => 
                           pipeline_stageD_offset_jump_sign_ext_24_port, A2 => 
                           n17328, A3 => n17315, ZN => n16533);
   U12231 : NAND3_X1 port map( A1 => 
                           pipeline_stageD_offset_jump_sign_ext_31_port, A2 => 
                           pipeline_stageD_offset_jump_sign_ext_24_port, A3 => 
                           n17315, ZN => n16545);
   U12232 : NAND3_X1 port map( A1 => 
                           pipeline_stageD_offset_jump_sign_ext_24_port, A2 => 
                           pipeline_stageD_offset_jump_sign_ext_31_port, A3 => 
                           pipeline_stageD_offset_jump_sign_ext_21_port, ZN => 
                           n16546);
   U12235 : NAND3_X1 port map( A1 => pipeline_RegDst_to_WB_0_port, A2 => n17326
                           , A3 => n17304, ZN => n16576);
   U12236 : NAND3_X1 port map( A1 => pipeline_RegDst_to_WB_1_port, A2 => n17314
                           , A3 => n17326, ZN => n16578);
   U12237 : NAND3_X1 port map( A1 => pipeline_RegDst_to_WB_0_port, A2 => 
                           pipeline_RegDst_to_WB_1_port, A3 => n17326, ZN => 
                           n16579);
   U12238 : NAND3_X1 port map( A1 => pipeline_RegDst_to_WB_2_port, A2 => n17314
                           , A3 => n17304, ZN => n16580);
   U12239 : NAND3_X1 port map( A1 => pipeline_RegDst_to_WB_2_port, A2 => 
                           pipeline_RegDst_to_WB_0_port, A3 => n17304, ZN => 
                           n16581);
   U12240 : NAND3_X1 port map( A1 => pipeline_RegDst_to_WB_2_port, A2 => 
                           pipeline_RegDst_to_WB_1_port, A3 => n17314, ZN => 
                           n16582);
   U12242 : NAND3_X1 port map( A1 => pipeline_RegDst_to_WB_0_port, A2 => 
                           pipeline_RegDst_to_WB_2_port, A3 => 
                           pipeline_RegDst_to_WB_1_port, ZN => n16583);
   U12244 : NAND3_X1 port map( A1 => n16657, A2 => n15432, A3 => n15430, ZN => 
                           n16652);
   U12245 : XOR2_X1 port map( A => n17381, B => n15553, Z => n16677);
   U12246 : XOR2_X1 port map( A => n17381, B => n15512, Z => n15521);
   U12247 : XOR2_X1 port map( A => n17381, B => n15474, Z => n16666);
   U12248 : XOR2_X1 port map( A => n17381, B => n15449, Z => n15459);
   U12249 : XOR2_X1 port map( A => n17381, B => n15346, Z => n15348);
   U12250 : XOR2_X1 port map( A => n17381, B => n15312, Z => n16629);
   U12251 : XOR2_X1 port map( A => n17381, B => n15285, Z => n16626);
   U12252 : XOR2_X1 port map( A => n17381, B => n15261, Z => n15263);
   U12253 : XOR2_X1 port map( A => n17381, B => n15224, Z => n15234);
   U12254 : XOR2_X1 port map( A => n17381, B => n15216, Z => n16612);
   U12255 : XOR2_X1 port map( A => n17381, B => n15202, Z => n15204);
   U12256 : XOR2_X1 port map( A => n17381, B => n15182, Z => n16611);
   U12257 : NAND3_X1 port map( A1 => n16789, A2 => n16790, A3 => n16791, ZN => 
                           n16785);
   U12258 : XOR2_X1 port map( A => n17645, B => 
                           pipeline_Reg2_Addr_to_exe_1_port, Z => n16791);
   U12259 : XOR2_X1 port map( A => n17646, B => 
                           pipeline_Reg2_Addr_to_exe_2_port, Z => n16790);
   U12261 : XOR2_X1 port map( A => pipeline_regDst_to_mem_0_port, B => 
                           pipeline_Reg1_Addr_to_exe_0_port, Z => n16809);
   getInstr : IRAM port map( ck => Clk, Rst => Rst, Addr(31) => 
                           addr_to_iram_31_port, Addr(30) => 
                           addr_to_iram_30_port, Addr(29) => 
                           addr_to_iram_29_port, Addr(28) => 
                           addr_to_iram_28_port, Addr(27) => 
                           addr_to_iram_27_port, Addr(26) => 
                           addr_to_iram_26_port, Addr(25) => 
                           addr_to_iram_25_port, Addr(24) => 
                           addr_to_iram_24_port, Addr(23) => 
                           addr_to_iram_23_port, Addr(22) => 
                           addr_to_iram_22_port, Addr(21) => 
                           addr_to_iram_21_port, Addr(20) => 
                           addr_to_iram_20_port, Addr(19) => 
                           addr_to_iram_19_port, Addr(18) => 
                           addr_to_iram_18_port, Addr(17) => 
                           addr_to_iram_17_port, Addr(16) => 
                           addr_to_iram_16_port, Addr(15) => 
                           addr_to_iram_15_port, Addr(14) => 
                           addr_to_iram_14_port, Addr(13) => 
                           addr_to_iram_13_port, Addr(12) => 
                           addr_to_iram_12_port, Addr(11) => 
                           addr_to_iram_11_port, Addr(10) => 
                           addr_to_iram_10_port, Addr(9) => addr_to_iram_9_port
                           , Addr(8) => addr_to_iram_8_port, Addr(7) => 
                           addr_to_iram_7_port, Addr(6) => addr_to_iram_6_port,
                           Addr(5) => addr_to_iram_5_port, Addr(4) => 
                           addr_to_iram_4_port, Addr(3) => addr_to_iram_3_port,
                           Addr(2) => addr_to_iram_2_port, Addr(1) => 
                           pipeline_stageF_PC_plus4_N8, Addr(0) => 
                           pipeline_stageF_PC_plus4_N7, Dout(31) => 
                           InstrFetched_31_port, Dout(30) => 
                           InstrFetched_30_port, Dout(29) => 
                           InstrFetched_29_port, Dout(28) => 
                           InstrFetched_28_port, Dout(27) => 
                           InstrFetched_27_port, Dout(26) => 
                           InstrFetched_26_port, Dout(25) => 
                           InstrFetched_25_port, Dout(24) => 
                           InstrFetched_24_port, Dout(23) => 
                           InstrFetched_23_port, Dout(22) => 
                           InstrFetched_22_port, Dout(21) => 
                           InstrFetched_21_port, Dout(20) => 
                           InstrFetched_20_port, Dout(19) => 
                           InstrFetched_19_port, Dout(18) => 
                           InstrFetched_18_port, Dout(17) => 
                           InstrFetched_17_port, Dout(16) => 
                           InstrFetched_16_port, Dout(15) => 
                           InstrFetched_15_port, Dout(14) => 
                           InstrFetched_14_port, Dout(13) => 
                           InstrFetched_13_port, Dout(12) => 
                           InstrFetched_12_port, Dout(11) => 
                           InstrFetched_11_port, Dout(10) => 
                           InstrFetched_10_port, Dout(9) => InstrFetched_9_port
                           , Dout(8) => InstrFetched_8_port, Dout(7) => 
                           InstrFetched_7_port, Dout(6) => InstrFetched_6_port,
                           Dout(5) => InstrFetched_5_port, Dout(4) => 
                           InstrFetched_4_port, Dout(3) => InstrFetched_3_port,
                           Dout(2) => InstrFetched_2_port, Dout(1) => 
                           InstrFetched_1_port, Dout(0) => InstrFetched_0_port)
                           ;
   pipeline_stageD_evaluate_jump_target_targetJump_out_adder_tri_30_inst : 
                           TBUF_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_N63, EN => Rst,
                           Z => pipeline_stageD_target_Jump_temp_30_port);
   pipeline_stageD_evaluate_jump_target_targetJump_out_adder_tri_19_inst : 
                           TBUF_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_N52, EN => Rst,
                           Z => pipeline_stageD_target_Jump_temp_19_port);
   pipeline_stageD_evaluate_jump_target_targetJump_out_adder_tri_21_inst : 
                           TBUF_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_N54, EN => Rst,
                           Z => pipeline_stageD_target_Jump_temp_21_port);
   pipeline_stageD_evaluate_jump_target_targetJump_out_adder_tri_22_inst : 
                           TBUF_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_N55, EN => Rst,
                           Z => pipeline_stageD_target_Jump_temp_22_port);
   U12260 : NAND3_X1 port map( A1 => n17314, A2 => n17326, A3 => n17304, ZN => 
                           n16586);
   pipeline_IFID_stage_PC_out_IFID_reg_0_inst : DFF_X1 port map( D => n3879, CK
                           => Clk, Q => pipeline_nextPC_IFID_DEC_0_port, QN => 
                           n17450);
   pipeline_IFID_stage_Instr_out_IFID_reg_24_inst : DFF_X1 port map( D => n3964
                           , CK => Clk, Q => 
                           pipeline_stageD_offset_jump_sign_ext_24_port, QN => 
                           n17384);
   pipeline_IFID_stage_Instr_out_IFID_reg_29_inst : DFF_X1 port map( D => n3959
                           , CK => Clk, Q => pipeline_inst_IFID_DEC_29_port, QN
                           => n17382);
   pipeline_IFID_stage_Instr_out_IFID_reg_5_inst : DFF_X1 port map( D => n3982,
                           CK => Clk, Q => 
                           pipeline_stageD_offset_to_jump_temp_5_port, QN => 
                           n17350);
   pipeline_IFID_stage_Instr_out_IFID_reg_25_inst : DFF_X1 port map( D => n3963
                           , CK => Clk, Q => 
                           pipeline_stageD_offset_jump_sign_ext_31_port, QN => 
                           n17328);
   pipeline_IDEX_Stage_EXE_controls_out_IDEX_reg_0_inst : DFF_X2 port map( D =>
                           pipeline_IDEX_Stage_N93, CK => Clk, Q => 
                           pipeline_EXE_controls_in_EXEcute_0_port, QN => 
                           n17327);
   pipeline_MEMWB_Stage_RegDst_Addr_out_MEMWB_reg_2_inst : DFF_X1 port map( D 
                           => pipeline_MEMWB_Stage_N45, CK => Clk, Q => 
                           pipeline_RegDst_to_WB_2_port, QN => n17326);
   pipeline_IFID_stage_Instr_out_IFID_reg_22_inst : DFF_X1 port map( D => n3966
                           , CK => Clk, Q => 
                           pipeline_stageD_offset_jump_sign_ext_22_port, QN => 
                           n17317);
   pipeline_IFID_stage_Instr_out_IFID_reg_21_inst : DFF_X1 port map( D => n3967
                           , CK => Clk, Q => 
                           pipeline_stageD_offset_jump_sign_ext_21_port, QN => 
                           n17315);
   pipeline_IFID_stage_Instr_out_IFID_reg_27_inst : DFF_X1 port map( D => n3961
                           , CK => Clk, Q => pipeline_inst_IFID_DEC_27_port, QN
                           => n17313);
   DataMem_Dataout_tri_31_inst : TBUF_X1 port map( A => DataMem_N2256, EN => 
                           DataMem_N0, Z => data_from_dram_31_port);
   DataMem_Dataout_tri_30_inst : TBUF_X1 port map( A => DataMem_N2259, EN => 
                           DataMem_N1, Z => data_from_dram_30_port);
   DataMem_Dataout_tri_29_inst : TBUF_X1 port map( A => DataMem_N2262, EN => 
                           DataMem_N2, Z => data_from_dram_29_port);
   DataMem_Dataout_tri_28_inst : TBUF_X1 port map( A => DataMem_N2265, EN => 
                           DataMem_N3, Z => data_from_dram_28_port);
   DataMem_Dataout_tri_27_inst : TBUF_X1 port map( A => DataMem_N2268, EN => 
                           DataMem_N4, Z => data_from_dram_27_port);
   DataMem_Dataout_tri_26_inst : TBUF_X1 port map( A => DataMem_N2271, EN => 
                           DataMem_N5, Z => data_from_dram_26_port);
   DataMem_Dataout_tri_25_inst : TBUF_X1 port map( A => DataMem_N2274, EN => 
                           DataMem_N6, Z => data_from_dram_25_port);
   DataMem_Dataout_tri_24_inst : TBUF_X1 port map( A => DataMem_N2277, EN => 
                           DataMem_N7, Z => data_from_dram_24_port);
   DataMem_Dataout_tri_23_inst : TBUF_X1 port map( A => DataMem_N2280, EN => 
                           DataMem_N8, Z => data_from_dram_23_port);
   DataMem_Dataout_tri_22_inst : TBUF_X1 port map( A => DataMem_N2283, EN => 
                           DataMem_N9, Z => data_from_dram_22_port);
   DataMem_Dataout_tri_21_inst : TBUF_X1 port map( A => DataMem_N2286, EN => 
                           DataMem_N10, Z => data_from_dram_21_port);
   DataMem_Dataout_tri_20_inst : TBUF_X1 port map( A => DataMem_N2289, EN => 
                           DataMem_N11, Z => data_from_dram_20_port);
   DataMem_Dataout_tri_19_inst : TBUF_X1 port map( A => DataMem_N2292, EN => 
                           DataMem_N12, Z => data_from_dram_19_port);
   DataMem_Dataout_tri_18_inst : TBUF_X1 port map( A => DataMem_N2295, EN => 
                           DataMem_N13, Z => data_from_dram_18_port);
   DataMem_Dataout_tri_17_inst : TBUF_X1 port map( A => DataMem_N2298, EN => 
                           DataMem_N14, Z => data_from_dram_17_port);
   DataMem_Dataout_tri_16_inst : TBUF_X1 port map( A => DataMem_N2301, EN => 
                           DataMem_N15, Z => data_from_dram_16_port);
   DataMem_Dataout_tri_15_inst : TBUF_X1 port map( A => DataMem_N2304, EN => 
                           DataMem_N16, Z => data_from_dram_15_port);
   DataMem_Dataout_tri_14_inst : TBUF_X1 port map( A => DataMem_N2307, EN => 
                           DataMem_N17, Z => data_from_dram_14_port);
   DataMem_Dataout_tri_13_inst : TBUF_X1 port map( A => DataMem_N2310, EN => 
                           DataMem_N18, Z => data_from_dram_13_port);
   DataMem_Dataout_tri_12_inst : TBUF_X1 port map( A => DataMem_N2313, EN => 
                           DataMem_N19, Z => data_from_dram_12_port);
   DataMem_Dataout_tri_11_inst : TBUF_X1 port map( A => DataMem_N2316, EN => 
                           DataMem_N20, Z => data_from_dram_11_port);
   DataMem_Dataout_tri_10_inst : TBUF_X1 port map( A => DataMem_N2319, EN => 
                           DataMem_N21, Z => data_from_dram_10_port);
   DataMem_Dataout_tri_9_inst : TBUF_X1 port map( A => DataMem_N2322, EN => 
                           DataMem_N22, Z => data_from_dram_9_port);
   DataMem_Dataout_tri_8_inst : TBUF_X1 port map( A => DataMem_N2325, EN => 
                           DataMem_N23, Z => data_from_dram_8_port);
   DataMem_Dataout_tri_7_inst : TBUF_X1 port map( A => DataMem_N2328, EN => 
                           DataMem_N24, Z => data_from_dram_7_port);
   DataMem_Dataout_tri_6_inst : TBUF_X1 port map( A => DataMem_N2331, EN => 
                           DataMem_N25, Z => data_from_dram_6_port);
   DataMem_Dataout_tri_5_inst : TBUF_X1 port map( A => DataMem_N2334, EN => 
                           DataMem_N26, Z => data_from_dram_5_port);
   DataMem_Dataout_tri_4_inst : TBUF_X1 port map( A => DataMem_N2337, EN => 
                           DataMem_N27, Z => data_from_dram_4_port);
   DataMem_Dataout_tri_3_inst : TBUF_X1 port map( A => DataMem_N2340, EN => 
                           DataMem_N28, Z => data_from_dram_3_port);
   DataMem_Dataout_tri_2_inst : TBUF_X1 port map( A => DataMem_N2343, EN => 
                           DataMem_N29, Z => data_from_dram_2_port);
   DataMem_Dataout_tri_1_inst : TBUF_X1 port map( A => DataMem_N2346, EN => 
                           DataMem_N30, Z => data_from_dram_1_port);
   DataMem_Dataout_tri_0_inst : TBUF_X1 port map( A => DataMem_N2349, EN => 
                           DataMem_N31, Z => data_from_dram_0_port);
   pipeline_stageD_evaluate_jump_target_targetJump_out_adder_tri_31_inst : 
                           TBUF_X1 port map( A => n415, EN => Rst, Z => 
                           pipeline_stageD_target_Jump_temp_31_port);
   pipeline_stageD_evaluate_jump_target_targetJump_out_adder_tri_1_inst : 
                           TBUF_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_N34, EN => Rst,
                           Z => pipeline_stageD_target_Jump_temp_1_port);
   pipeline_stageD_evaluate_jump_target_targetJump_out_adder_tri_0_inst : 
                           TBUF_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_N33, EN => Rst,
                           Z => pipeline_stageD_target_Jump_temp_0_port);
   pipeline_stageD_evaluate_jump_target_targetJump_out_adder_tri_11_inst : 
                           TBUF_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_N44, EN => Rst,
                           Z => pipeline_stageD_target_Jump_temp_11_port);
   pipeline_stageD_evaluate_jump_target_targetJump_out_adder_tri_12_inst : 
                           TBUF_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_N45, EN => Rst,
                           Z => pipeline_stageD_target_Jump_temp_12_port);
   pipeline_stageD_evaluate_jump_target_targetJump_out_adder_tri_8_inst : 
                           TBUF_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_N41, EN => Rst,
                           Z => pipeline_stageD_target_Jump_temp_8_port);
   pipeline_stageD_evaluate_jump_target_targetJump_out_adder_tri_7_inst : 
                           TBUF_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_N40, EN => Rst,
                           Z => pipeline_stageD_target_Jump_temp_7_port);
   pipeline_stageD_evaluate_jump_target_targetJump_out_adder_tri_6_inst : 
                           TBUF_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_N39, EN => Rst,
                           Z => pipeline_stageD_target_Jump_temp_6_port);
   pipeline_stageD_evaluate_jump_target_targetJump_out_adder_tri_15_inst : 
                           TBUF_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_N48, EN => Rst,
                           Z => pipeline_stageD_target_Jump_temp_15_port);
   pipeline_stageD_evaluate_jump_target_targetJump_out_adder_tri_13_inst : 
                           TBUF_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_N46, EN => Rst,
                           Z => pipeline_stageD_target_Jump_temp_13_port);
   pipeline_stageD_evaluate_jump_target_targetJump_out_adder_tri_9_inst : 
                           TBUF_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_N42, EN => Rst,
                           Z => pipeline_stageD_target_Jump_temp_9_port);
   pipeline_stageD_evaluate_jump_target_targetJump_out_adder_tri_5_inst : 
                           TBUF_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_N38, EN => Rst,
                           Z => pipeline_stageD_target_Jump_temp_5_port);
   pipeline_stageD_evaluate_jump_target_targetJump_out_adder_tri_3_inst : 
                           TBUF_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_N36, EN => Rst,
                           Z => pipeline_stageD_target_Jump_temp_3_port);
   pipeline_stageD_evaluate_jump_target_targetJump_out_adder_tri_14_inst : 
                           TBUF_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_N47, EN => Rst,
                           Z => pipeline_stageD_target_Jump_temp_14_port);
   pipeline_stageD_evaluate_jump_target_targetJump_out_adder_tri_2_inst : 
                           TBUF_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_N35, EN => Rst,
                           Z => pipeline_stageD_target_Jump_temp_2_port);
   pipeline_stageD_evaluate_jump_target_targetJump_out_adder_tri_10_inst : 
                           TBUF_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_N43, EN => Rst,
                           Z => pipeline_stageD_target_Jump_temp_10_port);
   pipeline_stageD_evaluate_jump_target_targetJump_out_adder_tri_4_inst : 
                           TBUF_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_N37, EN => Rst,
                           Z => pipeline_stageD_target_Jump_temp_4_port);
   pipeline_stageD_evaluate_jump_target_targetJump_out_adder_tri_29_inst : 
                           TBUF_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_N62, EN => Rst,
                           Z => pipeline_stageD_target_Jump_temp_29_port);
   pipeline_stageD_evaluate_jump_target_targetJump_out_adder_tri_17_inst : 
                           TBUF_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_N50, EN => Rst,
                           Z => pipeline_stageD_target_Jump_temp_17_port);
   pipeline_stageD_evaluate_jump_target_targetJump_out_adder_tri_16_inst : 
                           TBUF_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_N49, EN => Rst,
                           Z => pipeline_stageD_target_Jump_temp_16_port);
   pipeline_stageD_evaluate_jump_target_targetJump_out_adder_tri_23_inst : 
                           TBUF_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_N56, EN => Rst,
                           Z => pipeline_stageD_target_Jump_temp_23_port);
   pipeline_stageD_evaluate_jump_target_targetJump_out_adder_tri_26_inst : 
                           TBUF_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_N59, EN => Rst,
                           Z => pipeline_stageD_target_Jump_temp_26_port);
   pipeline_stageD_evaluate_jump_target_targetJump_out_adder_tri_28_inst : 
                           TBUF_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_N61, EN => Rst,
                           Z => pipeline_stageD_target_Jump_temp_28_port);
   pipeline_stageD_evaluate_jump_target_targetJump_out_adder_tri_27_inst : 
                           TBUF_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_N60, EN => Rst,
                           Z => pipeline_stageD_target_Jump_temp_27_port);
   pipeline_stageD_evaluate_jump_target_targetJump_out_adder_tri_25_inst : 
                           TBUF_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_N58, EN => Rst,
                           Z => pipeline_stageD_target_Jump_temp_25_port);
   pipeline_stageD_evaluate_jump_target_targetJump_out_adder_tri_20_inst : 
                           TBUF_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_N53, EN => Rst,
                           Z => pipeline_stageD_target_Jump_temp_20_port);
   pipeline_stageD_evaluate_jump_target_targetJump_out_adder_tri_18_inst : 
                           TBUF_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_N51, EN => Rst,
                           Z => pipeline_stageD_target_Jump_temp_18_port);
   pipeline_stageD_evaluate_jump_target_targetJump_out_adder_tri_24_inst : 
                           TBUF_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_N57, EN => Rst,
                           Z => pipeline_stageD_target_Jump_temp_24_port);
   pipeline_EXMEM_stage_RegDst_Addr_out_EXMEM_reg_1_inst : DFF_X1 port map( D 
                           => pipeline_EXMEM_stage_N72, CK => Clk, Q => 
                           pipeline_regDst_to_mem_1_port, QN => n17645);
   pipeline_EXMEM_stage_RegDst_Addr_out_EXMEM_reg_2_inst : DFF_X1 port map( D 
                           => pipeline_EXMEM_stage_N73, CK => Clk, Q => 
                           net214675, QN => n17646);
   pipeline_MEMWB_Stage_RegDst_Addr_out_MEMWB_reg_0_inst : DFF_X1 port map( D 
                           => pipeline_MEMWB_Stage_N43, CK => Clk, Q => 
                           pipeline_RegDst_to_WB_0_port, QN => n17314);
   U8434 : OAI21_X1 port map( B1 => n13967, B2 => n17317, A => n13969, ZN => 
                           pipeline_stageD_offset_to_jump_temp_22_port);
   U8437 : OAI21_X1 port map( B1 => n17349, B2 => n13967, A => n13969, ZN => 
                           pipeline_stageD_offset_to_jump_temp_19_port);
   U8438 : OAI21_X1 port map( B1 => n17408, B2 => n13967, A => n13969, ZN => 
                           pipeline_stageD_offset_to_jump_temp_18_port);
   U8439 : OAI21_X1 port map( B1 => n17329, B2 => n13967, A => n13969, ZN => 
                           pipeline_stageD_offset_to_jump_temp_17_port);
   U8440 : OAI21_X1 port map( B1 => n17316, B2 => n13967, A => n13969, ZN => 
                           pipeline_stageD_offset_to_jump_temp_16_port);
   U8436 : OAI21_X1 port map( B1 => n17407, B2 => n13967, A => n13969, ZN => 
                           pipeline_stageD_offset_to_jump_temp_20_port);
   U8435 : OAI21_X1 port map( B1 => n13967, B2 => n17315, A => n13969, ZN => 
                           pipeline_stageD_offset_to_jump_temp_21_port);
   U8433 : OAI21_X1 port map( B1 => n13967, B2 => n17383, A => n13969, ZN => 
                           pipeline_stageD_offset_to_jump_temp_23_port);
   U8432 : OAI21_X1 port map( B1 => n13967, B2 => n17384, A => n13969, ZN => 
                           pipeline_stageD_offset_to_jump_temp_24_port);
   U10941 : OAI22_X1 port map( A1 => pipeline_regDst_to_mem_0_port, A2 => 
                           n17315, B1 => n17646, B2 => 
                           pipeline_stageD_offset_jump_sign_ext_23_port, ZN => 
                           n16575);
   U10940 : AOI221_X1 port map( B1 => n17315, B2 => 
                           pipeline_regDst_to_mem_0_port, C1 => n17646, C2 => 
                           pipeline_stageD_offset_jump_sign_ext_23_port, A => 
                           n16575, ZN => n16574);
   U10937 : OAI221_X1 port map( B1 => pipeline_regDst_to_mem_1_port, B2 => 
                           n17317, C1 => n17645, C2 => 
                           pipeline_stageD_offset_jump_sign_ext_22_port, A => 
                           n16572, ZN => n16555);
   U10935 : AOI22_X1 port map( A1 => n17385, A2 => 
                           pipeline_stageD_offset_jump_sign_ext_24_port, B1 => 
                           n17314, B2 => 
                           pipeline_stageD_offset_jump_sign_ext_21_port, ZN => 
                           n16571);
   U10934 : OAI221_X1 port map( B1 => n17385, B2 => 
                           pipeline_stageD_offset_jump_sign_ext_24_port, C1 => 
                           n17314, C2 => 
                           pipeline_stageD_offset_jump_sign_ext_21_port, A => 
                           n16571, ZN => n16562);
   U10928 : NOR4_X1 port map( A1 => pipeline_Alu_Out_Addr_to_mem_19_port, A2 =>
                           pipeline_Alu_Out_Addr_to_mem_18_port, A3 => 
                           pipeline_Alu_Out_Addr_to_mem_20_port, A4 => 
                           pipeline_Alu_Out_Addr_to_mem_21_port, ZN => n16556);
   U10927 : NOR4_X1 port map( A1 => pipeline_Alu_Out_Addr_to_mem_25_port, A2 =>
                           pipeline_Alu_Out_Addr_to_mem_24_port, A3 => 
                           pipeline_Alu_Out_Addr_to_mem_23_port, A4 => 
                           pipeline_Alu_Out_Addr_to_mem_22_port, ZN => n16557);
   U10926 : NOR4_X1 port map( A1 => pipeline_Alu_Out_Addr_to_mem_13_port, A2 =>
                           pipeline_Alu_Out_Addr_to_mem_11_port, A3 => 
                           pipeline_Alu_Out_Addr_to_mem_10_port, A4 => 
                           pipeline_Alu_Out_Addr_to_mem_12_port, ZN => n16558);
   U10925 : NOR4_X1 port map( A1 => pipeline_Alu_Out_Addr_to_mem_14_port, A2 =>
                           pipeline_Alu_Out_Addr_to_mem_15_port, A3 => 
                           pipeline_Alu_Out_Addr_to_mem_17_port, A4 => 
                           pipeline_Alu_Out_Addr_to_mem_16_port, ZN => n16559);
   U10924 : NAND4_X1 port map( A1 => n16556, A2 => n16557, A3 => n16558, A4 => 
                           n16559, ZN => n15887);
   U10921 : NOR4_X1 port map( A1 => pipeline_Alu_Out_Addr_to_mem_0_port, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_2_port, A3 => 
                           pipeline_Alu_Out_Addr_to_mem_1_port, A4 => 
                           pipeline_Alu_Out_Addr_to_mem_3_port, ZN => n16550);
   U10920 : NOR4_X1 port map( A1 => pipeline_Alu_Out_Addr_to_mem_8_port, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_7_port, A3 => 
                           pipeline_Alu_Out_Addr_to_mem_6_port, A4 => 
                           pipeline_Alu_Out_Addr_to_mem_9_port, ZN => n16551);
   U10919 : NOR4_X1 port map( A1 => pipeline_Alu_Out_Addr_to_mem_31_port, A2 =>
                           pipeline_Alu_Out_Addr_to_mem_4_port, A3 => 
                           pipeline_Alu_Out_Addr_to_mem_5_port, A4 => 
                           pipeline_Alu_Out_Addr_to_mem_30_port, ZN => n16552);
   U10918 : NOR4_X1 port map( A1 => pipeline_Alu_Out_Addr_to_mem_26_port, A2 =>
                           pipeline_Alu_Out_Addr_to_mem_27_port, A3 => 
                           pipeline_Alu_Out_Addr_to_mem_28_port, A4 => 
                           pipeline_Alu_Out_Addr_to_mem_29_port, ZN => n16553);
   U10917 : NAND4_X1 port map( A1 => n16550, A2 => n16551, A3 => n16552, A4 => 
                           n16553, ZN => n15888);
   U10913 : AOI22_X1 port map( A1 => n17137, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_31_26_port, B1 => 
                           n17138, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_26_port, ZN => 
                           n16547);
   U10909 : AOI22_X1 port map( A1 => n17130, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_29_26_port, B1 => 
                           n17129, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_26_port, ZN => 
                           n16548);
   U10904 : AOI222_X1 port map( A1 => n17135, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_8_26_port, B1 => 
                           n17132, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_26_port, C1 => 
                           n17127, C2 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_26_port, ZN => 
                           n16549);
   U10900 : AOI22_X1 port map( A1 => n17143, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_27_26_port, B1 => 
                           n17145, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_26_port, ZN => 
                           n16541);
   U10897 : AOI22_X1 port map( A1 => n17146, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_23_26_port, B1 => 
                           n17147, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_26_port, ZN => 
                           n16542);
   U10894 : AOI22_X1 port map( A1 => n17148, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_21_26_port, B1 => 
                           n17131, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_26_port, ZN => 
                           n16543);
   U10891 : AOI22_X1 port map( A1 => n17128, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_19_26_port, B1 => 
                           n17134, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_26_port, ZN => 
                           n16544);
   U10890 : NAND4_X1 port map( A1 => n16541, A2 => n16542, A3 => n16543, A4 => 
                           n16544, ZN => n16520);
   U10887 : AOI22_X1 port map( A1 => n17141, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_17_26_port, B1 => 
                           n17341, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_26_port, ZN => 
                           n16535);
   U10884 : AOI22_X1 port map( A1 => n17388, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_9_26_port, B1 => 
                           n17139, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_2_26_port, ZN => 
                           n16536);
   U10881 : AOI22_X1 port map( A1 => n17136, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_12_26_port, B1 => 
                           n17389, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_11_26_port, ZN => 
                           n16537);
   U10878 : AOI22_X1 port map( A1 => n17140, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_14_26_port, B1 => 
                           n17390, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_26_port, ZN => 
                           n16538);
   U10877 : NAND4_X1 port map( A1 => n16535, A2 => n16536, A3 => n16537, A4 => 
                           n16538, ZN => n16521);
   U10874 : AOI22_X1 port map( A1 => n17133, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_26_port, B1 => 
                           n17392, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_4_26_port, ZN => 
                           n16523);
   U10871 : AOI22_X1 port map( A1 => n17334, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_26_port, B1 => 
                           n17144, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_26_port, ZN => 
                           n16524);
   U10868 : AOI22_X1 port map( A1 => n17338, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_6_26_port, B1 => 
                           n17142, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_26_port, ZN => 
                           n16525);
   U10865 : AOI22_X1 port map( A1 => n17336, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_26_port, B1 => 
                           n17391, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_26_port, ZN => 
                           n16526);
   U10864 : NAND4_X1 port map( A1 => n16523, A2 => n16524, A3 => n16525, A4 => 
                           n16526, ZN => n16522);
   U10863 : NOR4_X1 port map( A1 => n16519, A2 => n16520, A3 => n16521, A4 => 
                           n16522, ZN => n14893);
   U10862 : AOI22_X1 port map( A1 => n15940, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_31_25_port, B1 => 
                           n15941, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_25_port, ZN => 
                           n16516);
   U10861 : AOI22_X1 port map( A1 => n15938, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_29_25_port, B1 => 
                           n15939, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_25_port, ZN => 
                           n16517);
   U10860 : AOI222_X1 port map( A1 => n15935, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_8_25_port, B1 => 
                           n15936, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_25_port, C1 => 
                           n15937, C2 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_25_port, ZN => 
                           n16518);
   U10859 : AOI22_X1 port map( A1 => n15930, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_27_25_port, B1 => 
                           n15931, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_25_port, ZN => 
                           n16512);
   U10858 : AOI22_X1 port map( A1 => n15928, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_23_25_port, B1 => 
                           n15929, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_25_port, ZN => 
                           n16513);
   U10857 : AOI22_X1 port map( A1 => n15926, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_21_25_port, B1 => 
                           n15927, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_25_port, ZN => 
                           n16514);
   U10856 : AOI22_X1 port map( A1 => n15924, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_19_25_port, B1 => 
                           n15925, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_25_port, ZN => 
                           n16515);
   U10855 : NAND4_X1 port map( A1 => n16512, A2 => n16513, A3 => n16514, A4 => 
                           n16515, ZN => n16501);
   U10854 : AOI22_X1 port map( A1 => n15918, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_17_25_port, B1 => 
                           n17341, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_25_port, ZN => 
                           n16508);
   U10853 : AOI22_X1 port map( A1 => n17388, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_9_25_port, B1 => 
                           n15917, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_2_25_port, ZN => 
                           n16509);
   U10852 : AOI22_X1 port map( A1 => n15914, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_12_25_port, B1 => 
                           n17389, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_11_25_port, ZN => 
                           n16510);
   U10851 : AOI22_X1 port map( A1 => n15912, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_14_25_port, B1 => 
                           n17390, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_25_port, ZN => 
                           n16511);
   U10850 : NAND4_X1 port map( A1 => n16508, A2 => n16509, A3 => n16510, A4 => 
                           n16511, ZN => n16502);
   U10849 : AOI22_X1 port map( A1 => n15906, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_25_port, B1 => 
                           n17392, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_4_25_port, ZN => 
                           n16504);
   U10848 : AOI22_X1 port map( A1 => n17334, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_25_port, B1 => 
                           n15905, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_25_port, ZN => 
                           n16505);
   U10847 : AOI22_X1 port map( A1 => n17338, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_6_25_port, B1 => 
                           n15903, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_25_port, ZN => 
                           n16506);
   U10846 : AOI22_X1 port map( A1 => n17336, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_25_port, B1 => 
                           n17391, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_25_port, ZN => 
                           n16507);
   U10845 : NAND4_X1 port map( A1 => n16504, A2 => n16505, A3 => n16506, A4 => 
                           n16507, ZN => n16503);
   U10844 : NOR4_X1 port map( A1 => n16500, A2 => n16501, A3 => n16502, A4 => 
                           n16503, ZN => n14895);
   U10843 : AOI22_X1 port map( A1 => n17137, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_31_24_port, B1 => 
                           n17138, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_24_port, ZN => 
                           n16497);
   U10842 : AOI22_X1 port map( A1 => n17130, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_29_24_port, B1 => 
                           n17129, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_24_port, ZN => 
                           n16498);
   U10841 : AOI222_X1 port map( A1 => n17135, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_8_24_port, B1 => 
                           n17132, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_24_port, C1 => 
                           n17127, C2 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_24_port, ZN => 
                           n16499);
   U10840 : AOI22_X1 port map( A1 => n17143, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_27_24_port, B1 => 
                           n17145, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_24_port, ZN => 
                           n16493);
   U10839 : AOI22_X1 port map( A1 => n17146, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_23_24_port, B1 => 
                           n17147, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_24_port, ZN => 
                           n16494);
   U10838 : AOI22_X1 port map( A1 => n17148, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_21_24_port, B1 => 
                           n17131, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_24_port, ZN => 
                           n16495);
   U10837 : AOI22_X1 port map( A1 => n17128, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_19_24_port, B1 => 
                           n17134, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_24_port, ZN => 
                           n16496);
   U10836 : NAND4_X1 port map( A1 => n16493, A2 => n16494, A3 => n16495, A4 => 
                           n16496, ZN => n16482);
   U10835 : AOI22_X1 port map( A1 => n17141, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_17_24_port, B1 => 
                           n17341, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_24_port, ZN => 
                           n16489);
   U10834 : AOI22_X1 port map( A1 => n17388, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_9_24_port, B1 => 
                           n17139, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_2_24_port, ZN => 
                           n16490);
   U10833 : AOI22_X1 port map( A1 => n17136, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_12_24_port, B1 => 
                           n17389, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_11_24_port, ZN => 
                           n16491);
   U10832 : AOI22_X1 port map( A1 => n17140, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_14_24_port, B1 => 
                           n17390, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_24_port, ZN => 
                           n16492);
   U10831 : NAND4_X1 port map( A1 => n16489, A2 => n16490, A3 => n16491, A4 => 
                           n16492, ZN => n16483);
   U10830 : AOI22_X1 port map( A1 => n17133, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_24_port, B1 => 
                           n17392, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_4_24_port, ZN => 
                           n16485);
   U10829 : AOI22_X1 port map( A1 => n17334, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_24_port, B1 => 
                           n17144, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_24_port, ZN => 
                           n16486);
   U10828 : AOI22_X1 port map( A1 => n17338, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_6_24_port, B1 => 
                           n17142, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_24_port, ZN => 
                           n16487);
   U10827 : AOI22_X1 port map( A1 => n17336, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_24_port, B1 => 
                           n17391, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_24_port, ZN => 
                           n16488);
   U10826 : NAND4_X1 port map( A1 => n16485, A2 => n16486, A3 => n16487, A4 => 
                           n16488, ZN => n16484);
   U10825 : NOR4_X1 port map( A1 => n16481, A2 => n16482, A3 => n16483, A4 => 
                           n16484, ZN => n14897);
   U10824 : AOI22_X1 port map( A1 => n17137, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_31_23_port, B1 => 
                           n17138, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_23_port, ZN => 
                           n16478);
   U10823 : AOI22_X1 port map( A1 => n17130, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_29_23_port, B1 => 
                           n17129, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_23_port, ZN => 
                           n16479);
   U10822 : AOI222_X1 port map( A1 => n17135, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_8_23_port, B1 => 
                           n17132, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_23_port, C1 => 
                           n17127, C2 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_23_port, ZN => 
                           n16480);
   U10821 : AOI22_X1 port map( A1 => n17143, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_27_23_port, B1 => 
                           n17145, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_23_port, ZN => 
                           n16474);
   U10820 : AOI22_X1 port map( A1 => n17146, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_23_23_port, B1 => 
                           n17147, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_23_port, ZN => 
                           n16475);
   U10819 : AOI22_X1 port map( A1 => n17148, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_21_23_port, B1 => 
                           n17131, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_23_port, ZN => 
                           n16476);
   U10818 : AOI22_X1 port map( A1 => n17128, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_19_23_port, B1 => 
                           n17134, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_23_port, ZN => 
                           n16477);
   U10817 : NAND4_X1 port map( A1 => n16474, A2 => n16475, A3 => n16476, A4 => 
                           n16477, ZN => n16463);
   U10816 : AOI22_X1 port map( A1 => n17141, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_17_23_port, B1 => 
                           n17341, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_23_port, ZN => 
                           n16470);
   U10815 : AOI22_X1 port map( A1 => n17388, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_9_23_port, B1 => 
                           n17139, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_2_23_port, ZN => 
                           n16471);
   U10814 : AOI22_X1 port map( A1 => n17136, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_12_23_port, B1 => 
                           n17389, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_11_23_port, ZN => 
                           n16472);
   U10813 : AOI22_X1 port map( A1 => n17140, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_14_23_port, B1 => 
                           n17390, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_23_port, ZN => 
                           n16473);
   U10812 : NAND4_X1 port map( A1 => n16470, A2 => n16471, A3 => n16472, A4 => 
                           n16473, ZN => n16464);
   U10811 : AOI22_X1 port map( A1 => n17133, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_23_port, B1 => 
                           n17392, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_4_23_port, ZN => 
                           n16466);
   U10810 : AOI22_X1 port map( A1 => n17334, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_23_port, B1 => 
                           n17144, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_23_port, ZN => 
                           n16467);
   U10809 : AOI22_X1 port map( A1 => n17338, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_6_23_port, B1 => 
                           n17142, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_23_port, ZN => 
                           n16468);
   U10808 : AOI22_X1 port map( A1 => n17336, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_23_port, B1 => 
                           n17391, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_23_port, ZN => 
                           n16469);
   U10807 : NAND4_X1 port map( A1 => n16466, A2 => n16467, A3 => n16468, A4 => 
                           n16469, ZN => n16465);
   U10806 : NOR4_X1 port map( A1 => n16462, A2 => n16463, A3 => n16464, A4 => 
                           n16465, ZN => n14899);
   U10805 : NAND4_X1 port map( A1 => n14893, A2 => n14895, A3 => n14897, A4 => 
                           n14899, ZN => n15889);
   U10804 : AOI22_X1 port map( A1 => n17137, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_31_6_port, B1 => 
                           n17138, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_6_port, ZN => 
                           n16459);
   U10803 : AOI22_X1 port map( A1 => n17130, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_29_6_port, B1 => 
                           n17129, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_6_port, ZN => 
                           n16460);
   U10802 : AOI222_X1 port map( A1 => n17135, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_8_6_port, B1 => 
                           n17132, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_6_port, C1 => 
                           n17127, C2 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_6_port, ZN => 
                           n16461);
   U10801 : AOI22_X1 port map( A1 => n17143, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_27_6_port, B1 => 
                           n17145, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_6_port, ZN => 
                           n16455);
   U10800 : AOI22_X1 port map( A1 => n17146, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_23_6_port, B1 => 
                           n17147, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_6_port, ZN => 
                           n16456);
   U10799 : AOI22_X1 port map( A1 => n17148, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_21_6_port, B1 => 
                           n17131, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_6_port, ZN => 
                           n16457);
   U10798 : AOI22_X1 port map( A1 => n17128, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_19_6_port, B1 => 
                           n17134, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_6_port, ZN => 
                           n16458);
   U10797 : NAND4_X1 port map( A1 => n16455, A2 => n16456, A3 => n16457, A4 => 
                           n16458, ZN => n16444);
   U10796 : AOI22_X1 port map( A1 => n17141, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_17_6_port, B1 => 
                           n17342, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_6_port, ZN => 
                           n16451);
   U10795 : AOI22_X1 port map( A1 => n17388, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_9_6_port, B1 => 
                           n17139, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_2_6_port, ZN => 
                           n16452);
   U10794 : AOI22_X1 port map( A1 => n17136, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_12_6_port, B1 => 
                           n17389, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_11_6_port, ZN => 
                           n16453);
   U10793 : AOI22_X1 port map( A1 => n17140, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_14_6_port, B1 => 
                           n17390, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_6_port, ZN => 
                           n16454);
   U10792 : NAND4_X1 port map( A1 => n16451, A2 => n16452, A3 => n16453, A4 => 
                           n16454, ZN => n16445);
   U10791 : AOI22_X1 port map( A1 => n17133, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_6_port, B1 => 
                           n17392, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_4_6_port, ZN => 
                           n16447);
   U10790 : AOI22_X1 port map( A1 => n17335, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_6_port, B1 => 
                           n17144, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_6_port, ZN => 
                           n16448);
   U10789 : AOI22_X1 port map( A1 => n17339, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_6_6_port, B1 => 
                           n17142, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_6_port, ZN => 
                           n16449);
   U10788 : AOI22_X1 port map( A1 => n17337, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_6_port, B1 => 
                           n17391, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_6_port, ZN => 
                           n16450);
   U10787 : NAND4_X1 port map( A1 => n16447, A2 => n16448, A3 => n16449, A4 => 
                           n16450, ZN => n16446);
   U10786 : NOR4_X1 port map( A1 => n16443, A2 => n16444, A3 => n16445, A4 => 
                           n16446, ZN => n14933);
   U10785 : AOI22_X1 port map( A1 => n15940, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_31_5_port, B1 => 
                           n15941, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_5_port, ZN => 
                           n16440);
   U10784 : AOI22_X1 port map( A1 => n15938, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_29_5_port, B1 => 
                           n15939, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_5_port, ZN => 
                           n16441);
   U10783 : AOI222_X1 port map( A1 => n15935, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_8_5_port, B1 => 
                           n15936, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_5_port, C1 => 
                           n15937, C2 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_5_port, ZN => 
                           n16442);
   U10782 : AOI22_X1 port map( A1 => n15930, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_27_5_port, B1 => 
                           n15931, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_5_port, ZN => 
                           n16436);
   U10781 : AOI22_X1 port map( A1 => n15928, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_23_5_port, B1 => 
                           n15929, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_5_port, ZN => 
                           n16437);
   U10780 : AOI22_X1 port map( A1 => n15926, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_21_5_port, B1 => 
                           n15927, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_5_port, ZN => 
                           n16438);
   U10779 : AOI22_X1 port map( A1 => n15924, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_19_5_port, B1 => 
                           n15925, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_5_port, ZN => 
                           n16439);
   U10778 : NAND4_X1 port map( A1 => n16436, A2 => n16437, A3 => n16438, A4 => 
                           n16439, ZN => n16425);
   U10777 : AOI22_X1 port map( A1 => n15918, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_17_5_port, B1 => 
                           n17342, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_5_port, ZN => 
                           n16432);
   U10776 : AOI22_X1 port map( A1 => n17388, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_9_5_port, B1 => 
                           n15917, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_2_5_port, ZN => 
                           n16433);
   U10775 : AOI22_X1 port map( A1 => n15914, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_12_5_port, B1 => 
                           n17389, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_11_5_port, ZN => 
                           n16434);
   U10774 : AOI22_X1 port map( A1 => n15912, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_14_5_port, B1 => 
                           n17390, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_5_port, ZN => 
                           n16435);
   U10773 : NAND4_X1 port map( A1 => n16432, A2 => n16433, A3 => n16434, A4 => 
                           n16435, ZN => n16426);
   U10772 : AOI22_X1 port map( A1 => n15906, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_5_port, B1 => 
                           n17392, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_4_5_port, ZN => 
                           n16428);
   U10771 : AOI22_X1 port map( A1 => n17335, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_5_port, B1 => 
                           n15905, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_5_port, ZN => 
                           n16429);
   U10770 : AOI22_X1 port map( A1 => n17339, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_6_5_port, B1 => 
                           n15903, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_5_port, ZN => 
                           n16430);
   U10769 : AOI22_X1 port map( A1 => n17337, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_5_port, B1 => 
                           n17391, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_5_port, ZN => 
                           n16431);
   U10768 : NAND4_X1 port map( A1 => n16428, A2 => n16429, A3 => n16430, A4 => 
                           n16431, ZN => n16427);
   U10767 : NOR4_X1 port map( A1 => n16424, A2 => n16425, A3 => n16426, A4 => 
                           n16427, ZN => n14935);
   U10765 : AOI22_X1 port map( A1 => n15930, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_27_0_port, B1 => 
                           n15931, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_0_port, ZN => 
                           n16420);
   U10764 : AOI22_X1 port map( A1 => n15928, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_23_0_port, B1 => 
                           n15929, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_0_port, ZN => 
                           n16421);
   U10763 : AOI22_X1 port map( A1 => n15926, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_21_0_port, B1 => 
                           n15927, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_0_port, ZN => 
                           n16422);
   U10762 : AOI22_X1 port map( A1 => n15924, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_19_0_port, B1 => 
                           n15925, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_0_port, ZN => 
                           n16423);
   U10761 : NAND4_X1 port map( A1 => n16420, A2 => n16421, A3 => n16422, A4 => 
                           n16423, ZN => n16405);
   U10760 : AOI22_X1 port map( A1 => n15940, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_31_0_port, B1 => 
                           n15941, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_0_port, ZN => 
                           n16417);
   U10759 : AOI22_X1 port map( A1 => n15938, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_29_0_port, B1 => 
                           n15939, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_0_port, ZN => 
                           n16418);
   U10758 : AOI222_X1 port map( A1 => n15935, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_8_0_port, B1 => 
                           n15936, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_0_port, C1 => 
                           n15937, C2 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_0_port, ZN => 
                           n16419);
   U10757 : AOI22_X1 port map( A1 => n15906, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_0_port, B1 => 
                           n17392, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_4_0_port, ZN => 
                           n16413);
   U10756 : AOI22_X1 port map( A1 => n17335, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_0_port, B1 => 
                           n15905, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_0_port, ZN => 
                           n16414);
   U10755 : AOI22_X1 port map( A1 => n17339, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_6_0_port, B1 => 
                           n15903, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_0_port, ZN => 
                           n16415);
   U10754 : AOI22_X1 port map( A1 => n17337, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_0_port, B1 => 
                           n17391, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_0_port, ZN => 
                           n16416);
   U10753 : NAND4_X1 port map( A1 => n16413, A2 => n16414, A3 => n16415, A4 => 
                           n16416, ZN => n16407);
   U10752 : AOI22_X1 port map( A1 => n15918, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_17_0_port, B1 => 
                           n17342, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_0_port, ZN => 
                           n16409);
   U10751 : AOI22_X1 port map( A1 => n17388, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_9_0_port, B1 => 
                           n15917, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_2_0_port, ZN => 
                           n16410);
   U10750 : AOI22_X1 port map( A1 => n15914, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_12_0_port, B1 => 
                           n17389, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_11_0_port, ZN => 
                           n16411);
   U10749 : AOI22_X1 port map( A1 => n15912, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_14_0_port, B1 => 
                           n17390, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_0_port, ZN => 
                           n16412);
   U10748 : NAND4_X1 port map( A1 => n16409, A2 => n16410, A3 => n16411, A4 => 
                           n16412, ZN => n16408);
   U10747 : NOR4_X1 port map( A1 => n16405, A2 => n16406, A3 => n16407, A4 => 
                           n16408, ZN => n14945);
   U10745 : AOI22_X1 port map( A1 => n17143, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_27_31_port, B1 => 
                           n17145, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_31_port, ZN => 
                           n16401);
   U10744 : AOI22_X1 port map( A1 => n17146, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_23_31_port, B1 => 
                           n17147, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_31_port, ZN => 
                           n16402);
   U10743 : AOI22_X1 port map( A1 => n17148, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_21_31_port, B1 => 
                           n17131, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_31_port, ZN => 
                           n16403);
   U10742 : AOI22_X1 port map( A1 => n17128, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_19_31_port, B1 => 
                           n17134, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_31_port, ZN => 
                           n16404);
   U10741 : NAND4_X1 port map( A1 => n16401, A2 => n16402, A3 => n16403, A4 => 
                           n16404, ZN => n16386);
   U10740 : AOI22_X1 port map( A1 => n17137, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_31_31_port, B1 => 
                           n17138, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_31_port, ZN => 
                           n16398);
   U10739 : AOI22_X1 port map( A1 => n17130, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_29_31_port, B1 => 
                           n17129, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_31_port, ZN => 
                           n16399);
   U10738 : AOI222_X1 port map( A1 => n17135, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_8_31_port, B1 => 
                           n17132, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_31_port, C1 => 
                           n17127, C2 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_31_port, ZN => 
                           n16400);
   U10737 : AOI22_X1 port map( A1 => n17133, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_31_port, B1 => 
                           n15907, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_4_31_port, ZN => 
                           n16394);
   U10736 : AOI22_X1 port map( A1 => n17335, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_31_port, B1 => 
                           n17144, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_31_port, ZN => 
                           n16395);
   U10735 : AOI22_X1 port map( A1 => n17339, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_6_31_port, B1 => 
                           n17142, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_31_port, ZN => 
                           n16396);
   U10734 : AOI22_X1 port map( A1 => n17337, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_31_port, B1 => 
                           n15901, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_31_port, ZN => 
                           n16397);
   U10733 : NAND4_X1 port map( A1 => n16394, A2 => n16395, A3 => n16396, A4 => 
                           n16397, ZN => n16388);
   U10732 : AOI22_X1 port map( A1 => n17141, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_17_31_port, B1 => 
                           n17342, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_31_port, ZN => 
                           n16390);
   U10731 : AOI22_X1 port map( A1 => n15916, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_9_31_port, B1 => 
                           n17139, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_2_31_port, ZN => 
                           n16391);
   U10730 : AOI22_X1 port map( A1 => n17136, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_12_31_port, B1 => 
                           n15915, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_11_31_port, ZN => 
                           n16392);
   U10729 : AOI22_X1 port map( A1 => n17140, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_14_31_port, B1 => 
                           n15913, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_31_port, ZN => 
                           n16393);
   U10728 : NAND4_X1 port map( A1 => n16390, A2 => n16391, A3 => n16392, A4 => 
                           n16393, ZN => n16389);
   U10727 : NOR4_X1 port map( A1 => n16386, A2 => n16387, A3 => n16388, A4 => 
                           n16389, ZN => n14883);
   U10725 : AOI22_X1 port map( A1 => n17137, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_31_4_port, B1 => 
                           n17138, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_4_port, ZN => 
                           n16383);
   U10724 : AOI22_X1 port map( A1 => n17130, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_29_4_port, B1 => 
                           n17129, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_4_port, ZN => 
                           n16384);
   U10723 : AOI222_X1 port map( A1 => n17135, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_8_4_port, B1 => 
                           n17132, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_4_port, C1 => 
                           n17127, C2 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_4_port, ZN => 
                           n16385);
   U10722 : AOI22_X1 port map( A1 => n17143, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_27_4_port, B1 => 
                           n17145, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_4_port, ZN => 
                           n16379);
   U10721 : AOI22_X1 port map( A1 => n17146, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_23_4_port, B1 => 
                           n17147, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_4_port, ZN => 
                           n16380);
   U10720 : AOI22_X1 port map( A1 => n17148, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_21_4_port, B1 => 
                           n17131, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_4_port, ZN => 
                           n16381);
   U10719 : AOI22_X1 port map( A1 => n17128, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_19_4_port, B1 => 
                           n17134, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_4_port, ZN => 
                           n16382);
   U10718 : NAND4_X1 port map( A1 => n16379, A2 => n16380, A3 => n16381, A4 => 
                           n16382, ZN => n16368);
   U10717 : AOI22_X1 port map( A1 => n17141, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_17_4_port, B1 => 
                           n17342, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_4_port, ZN => 
                           n16375);
   U10716 : AOI22_X1 port map( A1 => n15916, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_9_4_port, B1 => 
                           n17139, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_2_4_port, ZN => 
                           n16376);
   U10715 : AOI22_X1 port map( A1 => n17136, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_12_4_port, B1 => 
                           n15915, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_11_4_port, ZN => 
                           n16377);
   U10714 : AOI22_X1 port map( A1 => n17140, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_14_4_port, B1 => 
                           n15913, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_4_port, ZN => 
                           n16378);
   U10713 : NAND4_X1 port map( A1 => n16375, A2 => n16376, A3 => n16377, A4 => 
                           n16378, ZN => n16369);
   U10712 : AOI22_X1 port map( A1 => n17133, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_4_port, B1 => 
                           n15907, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_4_4_port, ZN => 
                           n16371);
   U10711 : AOI22_X1 port map( A1 => n17335, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_4_port, B1 => 
                           n17144, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_4_port, ZN => 
                           n16372);
   U10710 : AOI22_X1 port map( A1 => n17339, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_6_4_port, B1 => 
                           n17142, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_4_port, ZN => 
                           n16373);
   U10709 : AOI22_X1 port map( A1 => n17337, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_4_port, B1 => 
                           n15901, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_4_port, ZN => 
                           n16374);
   U10708 : NAND4_X1 port map( A1 => n16371, A2 => n16372, A3 => n16373, A4 => 
                           n16374, ZN => n16370);
   U10707 : NOR4_X1 port map( A1 => n16367, A2 => n16368, A3 => n16369, A4 => 
                           n16370, ZN => n14937);
   U10706 : AOI22_X1 port map( A1 => n17137, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_31_3_port, B1 => 
                           n17138, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_3_port, ZN => 
                           n16364);
   U10705 : AOI22_X1 port map( A1 => n17130, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_29_3_port, B1 => 
                           n17129, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_3_port, ZN => 
                           n16365);
   U10704 : AOI222_X1 port map( A1 => n17135, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_8_3_port, B1 => 
                           n17132, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_3_port, C1 => 
                           n17127, C2 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_3_port, ZN => 
                           n16366);
   U10703 : AOI22_X1 port map( A1 => n17143, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_27_3_port, B1 => 
                           n17145, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_3_port, ZN => 
                           n16360);
   U10702 : AOI22_X1 port map( A1 => n17146, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_23_3_port, B1 => 
                           n17147, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_3_port, ZN => 
                           n16361);
   U10701 : AOI22_X1 port map( A1 => n17148, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_21_3_port, B1 => 
                           n17131, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_3_port, ZN => 
                           n16362);
   U10700 : AOI22_X1 port map( A1 => n17128, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_19_3_port, B1 => 
                           n17134, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_3_port, ZN => 
                           n16363);
   U10699 : NAND4_X1 port map( A1 => n16360, A2 => n16361, A3 => n16362, A4 => 
                           n16363, ZN => n16349);
   U10698 : AOI22_X1 port map( A1 => n17141, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_17_3_port, B1 => 
                           n17342, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_3_port, ZN => 
                           n16356);
   U10697 : AOI22_X1 port map( A1 => n15916, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_9_3_port, B1 => 
                           n17139, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_2_3_port, ZN => 
                           n16357);
   U10696 : AOI22_X1 port map( A1 => n17136, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_12_3_port, B1 => 
                           n15915, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_11_3_port, ZN => 
                           n16358);
   U10695 : AOI22_X1 port map( A1 => n17140, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_14_3_port, B1 => 
                           n15913, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_3_port, ZN => 
                           n16359);
   U10694 : NAND4_X1 port map( A1 => n16356, A2 => n16357, A3 => n16358, A4 => 
                           n16359, ZN => n16350);
   U10693 : AOI22_X1 port map( A1 => n17133, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_3_port, B1 => 
                           n15907, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_4_3_port, ZN => 
                           n16352);
   U10692 : AOI22_X1 port map( A1 => n17335, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_3_port, B1 => 
                           n17144, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_3_port, ZN => 
                           n16353);
   U10691 : AOI22_X1 port map( A1 => n17339, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_6_3_port, B1 => 
                           n17142, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_3_port, ZN => 
                           n16354);
   U10690 : AOI22_X1 port map( A1 => n17337, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_3_port, B1 => 
                           n15901, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_3_port, ZN => 
                           n16355);
   U10689 : NAND4_X1 port map( A1 => n16352, A2 => n16353, A3 => n16354, A4 => 
                           n16355, ZN => n16351);
   U10688 : NOR4_X1 port map( A1 => n16348, A2 => n16349, A3 => n16350, A4 => 
                           n16351, ZN => n14939);
   U10687 : AOI22_X1 port map( A1 => n17137, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_31_2_port, B1 => 
                           n17138, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_2_port, ZN => 
                           n16345);
   U10686 : AOI22_X1 port map( A1 => n17130, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_29_2_port, B1 => 
                           n17129, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_2_port, ZN => 
                           n16346);
   U10685 : AOI222_X1 port map( A1 => n17135, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_8_2_port, B1 => 
                           n17132, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_2_port, C1 => 
                           n17127, C2 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_2_port, ZN => 
                           n16347);
   U10684 : AOI22_X1 port map( A1 => n17143, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_27_2_port, B1 => 
                           n17145, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_2_port, ZN => 
                           n16341);
   U10683 : AOI22_X1 port map( A1 => n17146, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_23_2_port, B1 => 
                           n17147, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_2_port, ZN => 
                           n16342);
   U10682 : AOI22_X1 port map( A1 => n17148, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_21_2_port, B1 => 
                           n17131, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_2_port, ZN => 
                           n16343);
   U10681 : AOI22_X1 port map( A1 => n17128, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_19_2_port, B1 => 
                           n17134, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_2_port, ZN => 
                           n16344);
   U10680 : NAND4_X1 port map( A1 => n16341, A2 => n16342, A3 => n16343, A4 => 
                           n16344, ZN => n16330);
   U10888 : NOR2_X1 port map( A1 => n16527, A2 => n16539, ZN => n15919);
   U10679 : AOI22_X1 port map( A1 => n17141, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_17_2_port, B1 => 
                           n15919, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_2_port, ZN => 
                           n16337);
   U10678 : AOI22_X1 port map( A1 => n15916, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_9_2_port, B1 => 
                           n17139, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_2_2_port, ZN => 
                           n16338);
   U10677 : AOI22_X1 port map( A1 => n17136, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_12_2_port, B1 => 
                           n15915, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_11_2_port, ZN => 
                           n16339);
   U10676 : AOI22_X1 port map( A1 => n17140, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_14_2_port, B1 => 
                           n15913, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_2_port, ZN => 
                           n16340);
   U10675 : NAND4_X1 port map( A1 => n16337, A2 => n16338, A3 => n16339, A4 => 
                           n16340, ZN => n16331);
   U10674 : AOI22_X1 port map( A1 => n17133, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_2_port, B1 => 
                           n15907, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_4_2_port, ZN => 
                           n16333);
   U10873 : NOR2_X1 port map( A1 => n16533, A2 => n16532, ZN => n15904);
   U10673 : AOI22_X1 port map( A1 => n15904, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_2_port, B1 => 
                           n17144, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_2_port, ZN => 
                           n16334);
   U10870 : NOR2_X1 port map( A1 => n16530, A2 => n16531, ZN => n15902);
   U10672 : AOI22_X1 port map( A1 => n15902, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_6_2_port, B1 => 
                           n17142, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_2_port, ZN => 
                           n16335);
   U10671 : AOI22_X1 port map( A1 => n17345, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_2_port, B1 => 
                           n15901, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_2_port, ZN => 
                           n16336);
   U10670 : NAND4_X1 port map( A1 => n16333, A2 => n16334, A3 => n16335, A4 => 
                           n16336, ZN => n16332);
   U10669 : NOR4_X1 port map( A1 => n16329, A2 => n16330, A3 => n16331, A4 => 
                           n16332, ZN => n14941);
   U10668 : AOI22_X1 port map( A1 => n17137, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_31_1_port, B1 => 
                           n17138, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_1_port, ZN => 
                           n16326);
   U10667 : AOI22_X1 port map( A1 => n17130, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_29_1_port, B1 => 
                           n17129, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_1_port, ZN => 
                           n16327);
   U10666 : AOI222_X1 port map( A1 => n17135, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_8_1_port, B1 => 
                           n17132, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_1_port, C1 => 
                           n17127, C2 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_1_port, ZN => 
                           n16328);
   U10665 : AOI22_X1 port map( A1 => n17143, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_27_1_port, B1 => 
                           n17145, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_1_port, ZN => 
                           n16322);
   U10664 : AOI22_X1 port map( A1 => n17146, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_23_1_port, B1 => 
                           n17147, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_1_port, ZN => 
                           n16323);
   U10663 : AOI22_X1 port map( A1 => n17148, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_21_1_port, B1 => 
                           n17131, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_1_port, ZN => 
                           n16324);
   U10662 : AOI22_X1 port map( A1 => n17128, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_19_1_port, B1 => 
                           n17134, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_1_port, ZN => 
                           n16325);
   U10661 : NAND4_X1 port map( A1 => n16322, A2 => n16323, A3 => n16324, A4 => 
                           n16325, ZN => n16311);
   U10660 : AOI22_X1 port map( A1 => n17141, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_17_1_port, B1 => 
                           n15919, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_1_port, ZN => 
                           n16318);
   U10659 : AOI22_X1 port map( A1 => n15916, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_9_1_port, B1 => 
                           n17139, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_2_1_port, ZN => 
                           n16319);
   U10658 : AOI22_X1 port map( A1 => n17136, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_12_1_port, B1 => 
                           n15915, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_11_1_port, ZN => 
                           n16320);
   U10657 : AOI22_X1 port map( A1 => n17140, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_14_1_port, B1 => 
                           n15913, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_1_port, ZN => 
                           n16321);
   U10656 : NAND4_X1 port map( A1 => n16318, A2 => n16319, A3 => n16320, A4 => 
                           n16321, ZN => n16312);
   U10655 : AOI22_X1 port map( A1 => n17133, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_1_port, B1 => 
                           n15907, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_4_1_port, ZN => 
                           n16314);
   U10654 : AOI22_X1 port map( A1 => n15904, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_1_port, B1 => 
                           n17144, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_1_port, ZN => 
                           n16315);
   U10653 : AOI22_X1 port map( A1 => n15902, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_6_1_port, B1 => 
                           n17142, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_1_port, ZN => 
                           n16316);
   U10652 : AOI22_X1 port map( A1 => n17345, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_1_port, B1 => 
                           n15901, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_1_port, ZN => 
                           n16317);
   U10651 : NAND4_X1 port map( A1 => n16314, A2 => n16315, A3 => n16316, A4 => 
                           n16317, ZN => n16313);
   U10650 : NOR4_X1 port map( A1 => n16310, A2 => n16311, A3 => n16312, A4 => 
                           n16313, ZN => n14943);
   U10649 : NAND4_X1 port map( A1 => n14937, A2 => n14939, A3 => n14941, A4 => 
                           n14943, ZN => n16309);
   U10648 : NOR4_X1 port map( A1 => n15832, A2 => n15772, A3 => n15688, A4 => 
                           n16309, ZN => n15999);
   U10647 : AOI22_X1 port map( A1 => n17137, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_31_18_port, B1 => 
                           n17138, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_18_port, ZN => 
                           n16306);
   U10646 : AOI22_X1 port map( A1 => n17130, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_29_18_port, B1 => 
                           n17129, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_18_port, ZN => 
                           n16307);
   U10645 : AOI222_X1 port map( A1 => n17135, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_8_18_port, B1 => 
                           n17132, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_18_port, C1 => 
                           n17127, C2 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_18_port, ZN => 
                           n16308);
   U10644 : AOI22_X1 port map( A1 => n17143, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_27_18_port, B1 => 
                           n17145, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_18_port, ZN => 
                           n16302);
   U10643 : AOI22_X1 port map( A1 => n17146, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_23_18_port, B1 => 
                           n17147, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_18_port, ZN => 
                           n16303);
   U10642 : AOI22_X1 port map( A1 => n17148, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_21_18_port, B1 => 
                           n17131, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_18_port, ZN => 
                           n16304);
   U10641 : AOI22_X1 port map( A1 => n17128, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_19_18_port, B1 => 
                           n17134, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_18_port, ZN => 
                           n16305);
   U10640 : NAND4_X1 port map( A1 => n16302, A2 => n16303, A3 => n16304, A4 => 
                           n16305, ZN => n16291);
   U10639 : AOI22_X1 port map( A1 => n17141, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_17_18_port, B1 => 
                           n15919, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_18_port, ZN => 
                           n16298);
   U10638 : AOI22_X1 port map( A1 => n15916, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_9_18_port, B1 => 
                           n17139, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_2_18_port, ZN => 
                           n16299);
   U10637 : AOI22_X1 port map( A1 => n17136, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_12_18_port, B1 => 
                           n15915, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_11_18_port, ZN => 
                           n16300);
   U10636 : AOI22_X1 port map( A1 => n17140, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_14_18_port, B1 => 
                           n15913, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_18_port, ZN => 
                           n16301);
   U10635 : NAND4_X1 port map( A1 => n16298, A2 => n16299, A3 => n16300, A4 => 
                           n16301, ZN => n16292);
   U10634 : AOI22_X1 port map( A1 => n17133, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_18_port, B1 => 
                           n15907, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_4_18_port, ZN => 
                           n16294);
   U10633 : AOI22_X1 port map( A1 => n15904, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_18_port, B1 => 
                           n17144, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_18_port, ZN => 
                           n16295);
   U10632 : AOI22_X1 port map( A1 => n15902, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_6_18_port, B1 => 
                           n17142, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_18_port, ZN => 
                           n16296);
   U10631 : AOI22_X1 port map( A1 => n17345, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_18_port, B1 => 
                           n15901, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_18_port, ZN => 
                           n16297);
   U10630 : NAND4_X1 port map( A1 => n16294, A2 => n16295, A3 => n16296, A4 => 
                           n16297, ZN => n16293);
   U10629 : NOR4_X1 port map( A1 => n16290, A2 => n16291, A3 => n16292, A4 => 
                           n16293, ZN => n14909);
   U10628 : AOI22_X1 port map( A1 => n17137, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_31_17_port, B1 => 
                           n17138, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_17_port, ZN => 
                           n16287);
   U10627 : AOI22_X1 port map( A1 => n17130, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_29_17_port, B1 => 
                           n17129, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_17_port, ZN => 
                           n16288);
   U10626 : AOI222_X1 port map( A1 => n17135, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_8_17_port, B1 => 
                           n17132, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_17_port, C1 => 
                           n17127, C2 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_17_port, ZN => 
                           n16289);
   U10625 : AOI22_X1 port map( A1 => n17143, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_27_17_port, B1 => 
                           n17145, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_17_port, ZN => 
                           n16283);
   U10624 : AOI22_X1 port map( A1 => n17146, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_23_17_port, B1 => 
                           n17147, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_17_port, ZN => 
                           n16284);
   U10623 : AOI22_X1 port map( A1 => n17148, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_21_17_port, B1 => 
                           n17131, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_17_port, ZN => 
                           n16285);
   U10622 : AOI22_X1 port map( A1 => n17128, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_19_17_port, B1 => 
                           n17134, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_17_port, ZN => 
                           n16286);
   U10621 : NAND4_X1 port map( A1 => n16283, A2 => n16284, A3 => n16285, A4 => 
                           n16286, ZN => n16272);
   U10620 : AOI22_X1 port map( A1 => n17141, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_17_17_port, B1 => 
                           n17341, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_17_port, ZN => 
                           n16279);
   U10619 : AOI22_X1 port map( A1 => n17388, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_9_17_port, B1 => 
                           n17139, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_2_17_port, ZN => 
                           n16280);
   U10618 : AOI22_X1 port map( A1 => n17136, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_12_17_port, B1 => 
                           n17389, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_11_17_port, ZN => 
                           n16281);
   U10617 : AOI22_X1 port map( A1 => n17140, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_14_17_port, B1 => 
                           n17390, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_17_port, ZN => 
                           n16282);
   U10616 : NAND4_X1 port map( A1 => n16279, A2 => n16280, A3 => n16281, A4 => 
                           n16282, ZN => n16273);
   U10615 : AOI22_X1 port map( A1 => n17133, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_17_port, B1 => 
                           n17392, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_4_17_port, ZN => 
                           n16275);
   U10614 : AOI22_X1 port map( A1 => n17334, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_17_port, B1 => 
                           n17144, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_17_port, ZN => 
                           n16276);
   U10613 : AOI22_X1 port map( A1 => n17338, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_6_17_port, B1 => 
                           n17142, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_17_port, ZN => 
                           n16277);
   U10612 : AOI22_X1 port map( A1 => n17336, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_17_port, B1 => 
                           n17391, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_17_port, ZN => 
                           n16278);
   U10611 : NAND4_X1 port map( A1 => n16275, A2 => n16276, A3 => n16277, A4 => 
                           n16278, ZN => n16274);
   U10610 : NOR4_X1 port map( A1 => n16271, A2 => n16272, A3 => n16273, A4 => 
                           n16274, ZN => n14911);
   U10609 : AOI22_X1 port map( A1 => n15940, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_31_16_port, B1 => 
                           n15941, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_16_port, ZN => 
                           n16268);
   U10608 : AOI22_X1 port map( A1 => n15938, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_29_16_port, B1 => 
                           n15939, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_16_port, ZN => 
                           n16269);
   U10607 : AOI222_X1 port map( A1 => n15935, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_8_16_port, B1 => 
                           n15936, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_16_port, C1 => 
                           n15937, C2 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_16_port, ZN => 
                           n16270);
   U10606 : AOI22_X1 port map( A1 => n15930, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_27_16_port, B1 => 
                           n15931, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_16_port, ZN => 
                           n16264);
   U10605 : AOI22_X1 port map( A1 => n15928, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_23_16_port, B1 => 
                           n15929, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_16_port, ZN => 
                           n16265);
   U10604 : AOI22_X1 port map( A1 => n15926, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_21_16_port, B1 => 
                           n15927, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_16_port, ZN => 
                           n16266);
   U10603 : AOI22_X1 port map( A1 => n15924, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_19_16_port, B1 => 
                           n15925, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_16_port, ZN => 
                           n16267);
   U10602 : NAND4_X1 port map( A1 => n16264, A2 => n16265, A3 => n16266, A4 => 
                           n16267, ZN => n16253);
   U10601 : AOI22_X1 port map( A1 => n15918, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_17_16_port, B1 => 
                           n17342, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_16_port, ZN => 
                           n16260);
   U10600 : AOI22_X1 port map( A1 => n15916, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_9_16_port, B1 => 
                           n15917, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_2_16_port, ZN => 
                           n16261);
   U10599 : AOI22_X1 port map( A1 => n15914, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_12_16_port, B1 => 
                           n15915, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_11_16_port, ZN => 
                           n16262);
   U10598 : AOI22_X1 port map( A1 => n15912, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_14_16_port, B1 => 
                           n15913, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_16_port, ZN => 
                           n16263);
   U10597 : NAND4_X1 port map( A1 => n16260, A2 => n16261, A3 => n16262, A4 => 
                           n16263, ZN => n16254);
   U10596 : AOI22_X1 port map( A1 => n15906, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_16_port, B1 => 
                           n15907, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_4_16_port, ZN => 
                           n16256);
   U10595 : AOI22_X1 port map( A1 => n17335, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_16_port, B1 => 
                           n15905, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_16_port, ZN => 
                           n16257);
   U10594 : AOI22_X1 port map( A1 => n17339, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_6_16_port, B1 => 
                           n15903, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_16_port, ZN => 
                           n16258);
   U10593 : AOI22_X1 port map( A1 => n17337, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_16_port, B1 => 
                           n15901, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_16_port, ZN => 
                           n16259);
   U10592 : NAND4_X1 port map( A1 => n16256, A2 => n16257, A3 => n16258, A4 => 
                           n16259, ZN => n16255);
   U10591 : NOR4_X1 port map( A1 => n16252, A2 => n16253, A3 => n16254, A4 => 
                           n16255, ZN => n14913);
   U10590 : AOI22_X1 port map( A1 => n15940, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_31_15_port, B1 => 
                           n15941, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_15_port, ZN => 
                           n16249);
   U10589 : AOI22_X1 port map( A1 => n15938, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_29_15_port, B1 => 
                           n15939, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_15_port, ZN => 
                           n16250);
   U10588 : AOI222_X1 port map( A1 => n15935, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_8_15_port, B1 => 
                           n15936, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_15_port, C1 => 
                           n15937, C2 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_15_port, ZN => 
                           n16251);
   U10587 : AOI22_X1 port map( A1 => n15930, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_27_15_port, B1 => 
                           n15931, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_15_port, ZN => 
                           n16245);
   U10586 : AOI22_X1 port map( A1 => n15928, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_23_15_port, B1 => 
                           n15929, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_15_port, ZN => 
                           n16246);
   U10585 : AOI22_X1 port map( A1 => n15926, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_21_15_port, B1 => 
                           n15927, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_15_port, ZN => 
                           n16247);
   U10584 : AOI22_X1 port map( A1 => n15924, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_19_15_port, B1 => 
                           n15925, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_15_port, ZN => 
                           n16248);
   U10583 : NAND4_X1 port map( A1 => n16245, A2 => n16246, A3 => n16247, A4 => 
                           n16248, ZN => n16234);
   U10582 : AOI22_X1 port map( A1 => n15918, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_17_15_port, B1 => 
                           n17342, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_15_port, ZN => 
                           n16241);
   U10581 : AOI22_X1 port map( A1 => n15916, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_9_15_port, B1 => 
                           n15917, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_2_15_port, ZN => 
                           n16242);
   U10580 : AOI22_X1 port map( A1 => n15914, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_12_15_port, B1 => 
                           n15915, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_11_15_port, ZN => 
                           n16243);
   U10579 : AOI22_X1 port map( A1 => n15912, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_14_15_port, B1 => 
                           n15913, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_15_port, ZN => 
                           n16244);
   U10578 : NAND4_X1 port map( A1 => n16241, A2 => n16242, A3 => n16243, A4 => 
                           n16244, ZN => n16235);
   U10577 : AOI22_X1 port map( A1 => n15906, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_15_port, B1 => 
                           n15907, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_4_15_port, ZN => 
                           n16237);
   U10576 : AOI22_X1 port map( A1 => n17335, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_15_port, B1 => 
                           n15905, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_15_port, ZN => 
                           n16238);
   U10575 : AOI22_X1 port map( A1 => n17339, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_6_15_port, B1 => 
                           n15903, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_15_port, ZN => 
                           n16239);
   U10574 : AOI22_X1 port map( A1 => n17337, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_15_port, B1 => 
                           n15901, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_15_port, ZN => 
                           n16240);
   U10573 : NAND4_X1 port map( A1 => n16237, A2 => n16238, A3 => n16239, A4 => 
                           n16240, ZN => n16236);
   U10572 : NOR4_X1 port map( A1 => n16233, A2 => n16234, A3 => n16235, A4 => 
                           n16236, ZN => n14915);
   U10571 : NAND4_X1 port map( A1 => n14909, A2 => n14911, A3 => n14913, A4 => 
                           n14915, ZN => n16001);
   U10570 : AOI22_X1 port map( A1 => n17137, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_31_22_port, B1 => 
                           n17138, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_22_port, ZN => 
                           n16230);
   U10569 : AOI22_X1 port map( A1 => n17130, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_29_22_port, B1 => 
                           n17129, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_22_port, ZN => 
                           n16231);
   U10568 : AOI222_X1 port map( A1 => n17135, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_8_22_port, B1 => 
                           n17132, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_22_port, C1 => 
                           n17127, C2 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_22_port, ZN => 
                           n16232);
   U10567 : AOI22_X1 port map( A1 => n17143, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_27_22_port, B1 => 
                           n17145, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_22_port, ZN => 
                           n16226);
   U10566 : AOI22_X1 port map( A1 => n17146, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_23_22_port, B1 => 
                           n17147, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_22_port, ZN => 
                           n16227);
   U10565 : AOI22_X1 port map( A1 => n17148, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_21_22_port, B1 => 
                           n17131, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_22_port, ZN => 
                           n16228);
   U10564 : AOI22_X1 port map( A1 => n17128, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_19_22_port, B1 => 
                           n17134, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_22_port, ZN => 
                           n16229);
   U10563 : NAND4_X1 port map( A1 => n16226, A2 => n16227, A3 => n16228, A4 => 
                           n16229, ZN => n16215);
   U10562 : AOI22_X1 port map( A1 => n17141, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_17_22_port, B1 => 
                           n15919, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_22_port, ZN => 
                           n16222);
   U10561 : AOI22_X1 port map( A1 => n15916, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_9_22_port, B1 => 
                           n17139, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_2_22_port, ZN => 
                           n16223);
   U10560 : AOI22_X1 port map( A1 => n17136, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_12_22_port, B1 => 
                           n15915, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_11_22_port, ZN => 
                           n16224);
   U10559 : AOI22_X1 port map( A1 => n17140, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_14_22_port, B1 => 
                           n15913, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_22_port, ZN => 
                           n16225);
   U10558 : NAND4_X1 port map( A1 => n16222, A2 => n16223, A3 => n16224, A4 => 
                           n16225, ZN => n16216);
   U10557 : AOI22_X1 port map( A1 => n17133, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_22_port, B1 => 
                           n15907, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_4_22_port, ZN => 
                           n16218);
   U10556 : AOI22_X1 port map( A1 => n15904, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_22_port, B1 => 
                           n17144, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_22_port, ZN => 
                           n16219);
   U10555 : AOI22_X1 port map( A1 => n15902, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_6_22_port, B1 => 
                           n17142, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_22_port, ZN => 
                           n16220);
   U10554 : AOI22_X1 port map( A1 => n17345, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_22_port, B1 => 
                           n15901, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_22_port, ZN => 
                           n16221);
   U10553 : NAND4_X1 port map( A1 => n16218, A2 => n16219, A3 => n16220, A4 => 
                           n16221, ZN => n16217);
   U10552 : NOR4_X1 port map( A1 => n16214, A2 => n16215, A3 => n16216, A4 => 
                           n16217, ZN => n14901);
   U10551 : AOI22_X1 port map( A1 => n17137, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_31_21_port, B1 => 
                           n17138, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_21_port, ZN => 
                           n16211);
   U10550 : AOI22_X1 port map( A1 => n17130, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_29_21_port, B1 => 
                           n17129, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_21_port, ZN => 
                           n16212);
   U10549 : AOI222_X1 port map( A1 => n17135, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_8_21_port, B1 => 
                           n17132, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_21_port, C1 => 
                           n17127, C2 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_21_port, ZN => 
                           n16213);
   U10548 : AOI22_X1 port map( A1 => n17143, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_27_21_port, B1 => 
                           n17145, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_21_port, ZN => 
                           n16207);
   U10547 : AOI22_X1 port map( A1 => n17146, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_23_21_port, B1 => 
                           n17147, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_21_port, ZN => 
                           n16208);
   U10546 : AOI22_X1 port map( A1 => n17148, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_21_21_port, B1 => 
                           n17131, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_21_port, ZN => 
                           n16209);
   U10545 : AOI22_X1 port map( A1 => n17128, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_19_21_port, B1 => 
                           n17134, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_21_port, ZN => 
                           n16210);
   U10544 : NAND4_X1 port map( A1 => n16207, A2 => n16208, A3 => n16209, A4 => 
                           n16210, ZN => n16196);
   U10543 : AOI22_X1 port map( A1 => n17141, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_17_21_port, B1 => 
                           n15919, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_21_port, ZN => 
                           n16203);
   U10542 : AOI22_X1 port map( A1 => n15916, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_9_21_port, B1 => 
                           n17139, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_2_21_port, ZN => 
                           n16204);
   U10541 : AOI22_X1 port map( A1 => n17136, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_12_21_port, B1 => 
                           n15915, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_11_21_port, ZN => 
                           n16205);
   U10540 : AOI22_X1 port map( A1 => n17140, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_14_21_port, B1 => 
                           n15913, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_21_port, ZN => 
                           n16206);
   U10539 : NAND4_X1 port map( A1 => n16203, A2 => n16204, A3 => n16205, A4 => 
                           n16206, ZN => n16197);
   U10538 : AOI22_X1 port map( A1 => n17133, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_21_port, B1 => 
                           n15907, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_4_21_port, ZN => 
                           n16199);
   U10537 : AOI22_X1 port map( A1 => n15904, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_21_port, B1 => 
                           n17144, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_21_port, ZN => 
                           n16200);
   U10536 : AOI22_X1 port map( A1 => n15902, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_6_21_port, B1 => 
                           n17142, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_21_port, ZN => 
                           n16201);
   U10535 : AOI22_X1 port map( A1 => n17345, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_21_port, B1 => 
                           n15901, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_21_port, ZN => 
                           n16202);
   U10534 : NAND4_X1 port map( A1 => n16199, A2 => n16200, A3 => n16201, A4 => 
                           n16202, ZN => n16198);
   U10533 : NOR4_X1 port map( A1 => n16195, A2 => n16196, A3 => n16197, A4 => 
                           n16198, ZN => n14903);
   U10532 : AOI22_X1 port map( A1 => n17137, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_31_20_port, B1 => 
                           n17138, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_20_port, ZN => 
                           n16192);
   U10531 : AOI22_X1 port map( A1 => n17130, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_29_20_port, B1 => 
                           n17129, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_20_port, ZN => 
                           n16193);
   U10530 : AOI222_X1 port map( A1 => n17135, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_8_20_port, B1 => 
                           n17132, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_20_port, C1 => 
                           n17127, C2 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_20_port, ZN => 
                           n16194);
   U10529 : AOI22_X1 port map( A1 => n17143, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_27_20_port, B1 => 
                           n17145, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_20_port, ZN => 
                           n16188);
   U10528 : AOI22_X1 port map( A1 => n17146, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_23_20_port, B1 => 
                           n17147, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_20_port, ZN => 
                           n16189);
   U10527 : AOI22_X1 port map( A1 => n17148, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_21_20_port, B1 => 
                           n17131, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_20_port, ZN => 
                           n16190);
   U10526 : AOI22_X1 port map( A1 => n17128, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_19_20_port, B1 => 
                           n17134, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_20_port, ZN => 
                           n16191);
   U10525 : NAND4_X1 port map( A1 => n16188, A2 => n16189, A3 => n16190, A4 => 
                           n16191, ZN => n16177);
   U10524 : AOI22_X1 port map( A1 => n17141, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_17_20_port, B1 => 
                           n15919, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_20_port, ZN => 
                           n16184);
   U10523 : AOI22_X1 port map( A1 => n15916, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_9_20_port, B1 => 
                           n17139, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_2_20_port, ZN => 
                           n16185);
   U10522 : AOI22_X1 port map( A1 => n17136, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_12_20_port, B1 => 
                           n15915, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_11_20_port, ZN => 
                           n16186);
   U10521 : AOI22_X1 port map( A1 => n17140, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_14_20_port, B1 => 
                           n15913, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_20_port, ZN => 
                           n16187);
   U10520 : NAND4_X1 port map( A1 => n16184, A2 => n16185, A3 => n16186, A4 => 
                           n16187, ZN => n16178);
   U10519 : AOI22_X1 port map( A1 => n17133, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_20_port, B1 => 
                           n15907, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_4_20_port, ZN => 
                           n16180);
   U10518 : AOI22_X1 port map( A1 => n15904, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_20_port, B1 => 
                           n17144, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_20_port, ZN => 
                           n16181);
   U10517 : AOI22_X1 port map( A1 => n15902, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_6_20_port, B1 => 
                           n17142, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_20_port, ZN => 
                           n16182);
   U10516 : AOI22_X1 port map( A1 => n17345, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_20_port, B1 => 
                           n15901, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_20_port, ZN => 
                           n16183);
   U10515 : NAND4_X1 port map( A1 => n16180, A2 => n16181, A3 => n16182, A4 => 
                           n16183, ZN => n16179);
   U10514 : NOR4_X1 port map( A1 => n16176, A2 => n16177, A3 => n16178, A4 => 
                           n16179, ZN => n14905);
   U10513 : AOI22_X1 port map( A1 => n15940, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_31_19_port, B1 => 
                           n15941, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_19_port, ZN => 
                           n16173);
   U10512 : AOI22_X1 port map( A1 => n15938, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_29_19_port, B1 => 
                           n15939, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_19_port, ZN => 
                           n16174);
   U10511 : AOI222_X1 port map( A1 => n15935, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_8_19_port, B1 => 
                           n15936, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_19_port, C1 => 
                           n15937, C2 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_19_port, ZN => 
                           n16175);
   U10510 : AOI22_X1 port map( A1 => n15930, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_27_19_port, B1 => 
                           n15931, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_19_port, ZN => 
                           n16169);
   U10509 : AOI22_X1 port map( A1 => n15928, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_23_19_port, B1 => 
                           n15929, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_19_port, ZN => 
                           n16170);
   U10508 : AOI22_X1 port map( A1 => n15926, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_21_19_port, B1 => 
                           n15927, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_19_port, ZN => 
                           n16171);
   U10507 : AOI22_X1 port map( A1 => n15924, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_19_19_port, B1 => 
                           n15925, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_19_port, ZN => 
                           n16172);
   U10506 : NAND4_X1 port map( A1 => n16169, A2 => n16170, A3 => n16171, A4 => 
                           n16172, ZN => n16158);
   U10505 : AOI22_X1 port map( A1 => n15918, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_17_19_port, B1 => 
                           n15919, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_19_port, ZN => 
                           n16165);
   U10504 : AOI22_X1 port map( A1 => n15916, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_9_19_port, B1 => 
                           n15917, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_2_19_port, ZN => 
                           n16166);
   U10503 : AOI22_X1 port map( A1 => n15914, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_12_19_port, B1 => 
                           n15915, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_11_19_port, ZN => 
                           n16167);
   U10502 : AOI22_X1 port map( A1 => n15912, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_14_19_port, B1 => 
                           n15913, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_19_port, ZN => 
                           n16168);
   U10501 : NAND4_X1 port map( A1 => n16165, A2 => n16166, A3 => n16167, A4 => 
                           n16168, ZN => n16159);
   U10500 : AOI22_X1 port map( A1 => n15906, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_19_port, B1 => 
                           n15907, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_4_19_port, ZN => 
                           n16161);
   U10499 : AOI22_X1 port map( A1 => n15904, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_19_port, B1 => 
                           n15905, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_19_port, ZN => 
                           n16162);
   U10498 : AOI22_X1 port map( A1 => n15902, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_6_19_port, B1 => 
                           n15903, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_19_port, ZN => 
                           n16163);
   U10497 : AOI22_X1 port map( A1 => n17345, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_19_port, B1 => 
                           n15901, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_19_port, ZN => 
                           n16164);
   U10496 : NAND4_X1 port map( A1 => n16161, A2 => n16162, A3 => n16163, A4 => 
                           n16164, ZN => n16160);
   U10495 : NOR4_X1 port map( A1 => n16157, A2 => n16158, A3 => n16159, A4 => 
                           n16160, ZN => n14907);
   U10494 : NAND4_X1 port map( A1 => n14901, A2 => n14903, A3 => n14905, A4 => 
                           n14907, ZN => n16002);
   U10493 : AOI22_X1 port map( A1 => n17137, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_31_10_port, B1 => 
                           n17138, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_10_port, ZN => 
                           n16154);
   U10492 : AOI22_X1 port map( A1 => n17130, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_29_10_port, B1 => 
                           n17129, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_10_port, ZN => 
                           n16155);
   U10491 : AOI222_X1 port map( A1 => n17135, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_8_10_port, B1 => 
                           n17132, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_10_port, C1 => 
                           n17127, C2 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_10_port, ZN => 
                           n16156);
   U10490 : AOI22_X1 port map( A1 => n17143, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_27_10_port, B1 => 
                           n17145, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_10_port, ZN => 
                           n16150);
   U10489 : AOI22_X1 port map( A1 => n17146, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_23_10_port, B1 => 
                           n17147, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_10_port, ZN => 
                           n16151);
   U10488 : AOI22_X1 port map( A1 => n17148, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_21_10_port, B1 => 
                           n17131, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_10_port, ZN => 
                           n16152);
   U10487 : AOI22_X1 port map( A1 => n17128, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_19_10_port, B1 => 
                           n17134, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_10_port, ZN => 
                           n16153);
   U10486 : NAND4_X1 port map( A1 => n16150, A2 => n16151, A3 => n16152, A4 => 
                           n16153, ZN => n16139);
   U10485 : AOI22_X1 port map( A1 => n17141, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_17_10_port, B1 => 
                           n15919, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_10_port, ZN => 
                           n16146);
   U10484 : AOI22_X1 port map( A1 => n15916, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_9_10_port, B1 => 
                           n17139, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_2_10_port, ZN => 
                           n16147);
   U10483 : AOI22_X1 port map( A1 => n17136, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_12_10_port, B1 => 
                           n15915, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_11_10_port, ZN => 
                           n16148);
   U10482 : AOI22_X1 port map( A1 => n17140, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_14_10_port, B1 => 
                           n15913, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_10_port, ZN => 
                           n16149);
   U10481 : NAND4_X1 port map( A1 => n16146, A2 => n16147, A3 => n16148, A4 => 
                           n16149, ZN => n16140);
   U10480 : AOI22_X1 port map( A1 => n17133, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_10_port, B1 => 
                           n15907, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_4_10_port, ZN => 
                           n16142);
   U10479 : AOI22_X1 port map( A1 => n15904, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_10_port, B1 => 
                           n17144, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_10_port, ZN => 
                           n16143);
   U10478 : AOI22_X1 port map( A1 => n15902, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_6_10_port, B1 => 
                           n17142, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_10_port, ZN => 
                           n16144);
   U10477 : AOI22_X1 port map( A1 => n17345, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_10_port, B1 => 
                           n15901, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_10_port, ZN => 
                           n16145);
   U10476 : NAND4_X1 port map( A1 => n16142, A2 => n16143, A3 => n16144, A4 => 
                           n16145, ZN => n16141);
   U10475 : NOR4_X1 port map( A1 => n16138, A2 => n16139, A3 => n16140, A4 => 
                           n16141, ZN => n14925);
   U10474 : AOI22_X1 port map( A1 => n17137, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_31_9_port, B1 => 
                           n17138, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_9_port, ZN => 
                           n16135);
   U10473 : AOI22_X1 port map( A1 => n17130, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_29_9_port, B1 => 
                           n17129, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_9_port, ZN => 
                           n16136);
   U10472 : AOI222_X1 port map( A1 => n17135, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_8_9_port, B1 => 
                           n17132, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_9_port, C1 => 
                           n17127, C2 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_9_port, ZN => 
                           n16137);
   U10471 : AOI22_X1 port map( A1 => n17143, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_27_9_port, B1 => 
                           n17145, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_9_port, ZN => 
                           n16131);
   U10470 : AOI22_X1 port map( A1 => n17146, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_23_9_port, B1 => 
                           n17147, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_9_port, ZN => 
                           n16132);
   U10469 : AOI22_X1 port map( A1 => n17148, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_21_9_port, B1 => 
                           n17131, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_9_port, ZN => 
                           n16133);
   U10468 : AOI22_X1 port map( A1 => n17128, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_19_9_port, B1 => 
                           n17134, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_9_port, ZN => 
                           n16134);
   U10467 : NAND4_X1 port map( A1 => n16131, A2 => n16132, A3 => n16133, A4 => 
                           n16134, ZN => n16120);
   U10466 : AOI22_X1 port map( A1 => n17141, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_17_9_port, B1 => 
                           n17341, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_9_port, ZN => 
                           n16127);
   U10465 : AOI22_X1 port map( A1 => n17388, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_9_9_port, B1 => 
                           n17139, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_2_9_port, ZN => 
                           n16128);
   U10464 : AOI22_X1 port map( A1 => n17136, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_12_9_port, B1 => 
                           n17389, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_11_9_port, ZN => 
                           n16129);
   U10463 : AOI22_X1 port map( A1 => n17140, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_14_9_port, B1 => 
                           n17390, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_9_port, ZN => 
                           n16130);
   U10462 : NAND4_X1 port map( A1 => n16127, A2 => n16128, A3 => n16129, A4 => 
                           n16130, ZN => n16121);
   U10461 : AOI22_X1 port map( A1 => n17133, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_9_port, B1 => 
                           n17392, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_4_9_port, ZN => 
                           n16123);
   U10460 : AOI22_X1 port map( A1 => n17334, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_9_port, B1 => 
                           n17144, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_9_port, ZN => 
                           n16124);
   U10459 : AOI22_X1 port map( A1 => n17338, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_6_9_port, B1 => 
                           n17142, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_9_port, ZN => 
                           n16125);
   U10458 : AOI22_X1 port map( A1 => n17336, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_9_port, B1 => 
                           n17391, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_9_port, ZN => 
                           n16126);
   U10457 : NAND4_X1 port map( A1 => n16123, A2 => n16124, A3 => n16125, A4 => 
                           n16126, ZN => n16122);
   U10456 : NOR4_X1 port map( A1 => n16119, A2 => n16120, A3 => n16121, A4 => 
                           n16122, ZN => n14927);
   U10455 : AOI22_X1 port map( A1 => n17137, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_31_8_port, B1 => 
                           n17138, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_8_port, ZN => 
                           n16116);
   U10454 : AOI22_X1 port map( A1 => n17130, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_29_8_port, B1 => 
                           n17129, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_8_port, ZN => 
                           n16117);
   U10453 : AOI222_X1 port map( A1 => n17135, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_8_8_port, B1 => 
                           n17132, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_8_port, C1 => 
                           n17127, C2 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_8_port, ZN => 
                           n16118);
   U10452 : AOI22_X1 port map( A1 => n17143, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_27_8_port, B1 => 
                           n17145, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_8_port, ZN => 
                           n16112);
   U10451 : AOI22_X1 port map( A1 => n17146, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_23_8_port, B1 => 
                           n17147, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_8_port, ZN => 
                           n16113);
   U10450 : AOI22_X1 port map( A1 => n17148, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_21_8_port, B1 => 
                           n17131, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_8_port, ZN => 
                           n16114);
   U10449 : AOI22_X1 port map( A1 => n17128, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_19_8_port, B1 => 
                           n17134, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_8_port, ZN => 
                           n16115);
   U10448 : NAND4_X1 port map( A1 => n16112, A2 => n16113, A3 => n16114, A4 => 
                           n16115, ZN => n16101);
   U10447 : AOI22_X1 port map( A1 => n17141, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_17_8_port, B1 => 
                           n17341, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_8_port, ZN => 
                           n16108);
   U10446 : AOI22_X1 port map( A1 => n17388, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_9_8_port, B1 => 
                           n17139, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_2_8_port, ZN => 
                           n16109);
   U10445 : AOI22_X1 port map( A1 => n17136, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_12_8_port, B1 => 
                           n17389, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_11_8_port, ZN => 
                           n16110);
   U10444 : AOI22_X1 port map( A1 => n17140, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_14_8_port, B1 => 
                           n17390, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_8_port, ZN => 
                           n16111);
   U10443 : NAND4_X1 port map( A1 => n16108, A2 => n16109, A3 => n16110, A4 => 
                           n16111, ZN => n16102);
   U10442 : AOI22_X1 port map( A1 => n17133, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_8_port, B1 => 
                           n17392, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_4_8_port, ZN => 
                           n16104);
   U10441 : AOI22_X1 port map( A1 => n17334, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_8_port, B1 => 
                           n17144, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_8_port, ZN => 
                           n16105);
   U10440 : AOI22_X1 port map( A1 => n17338, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_6_8_port, B1 => 
                           n17142, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_8_port, ZN => 
                           n16106);
   U10439 : AOI22_X1 port map( A1 => n17336, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_8_port, B1 => 
                           n17391, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_8_port, ZN => 
                           n16107);
   U10438 : NAND4_X1 port map( A1 => n16104, A2 => n16105, A3 => n16106, A4 => 
                           n16107, ZN => n16103);
   U10437 : NOR4_X1 port map( A1 => n16100, A2 => n16101, A3 => n16102, A4 => 
                           n16103, ZN => n14929);
   U10436 : AOI22_X1 port map( A1 => n17137, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_31_7_port, B1 => 
                           n17138, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_7_port, ZN => 
                           n16097);
   U10435 : AOI22_X1 port map( A1 => n17130, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_29_7_port, B1 => 
                           n17129, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_7_port, ZN => 
                           n16098);
   U10434 : AOI222_X1 port map( A1 => n17135, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_8_7_port, B1 => 
                           n17132, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_7_port, C1 => 
                           n17127, C2 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_7_port, ZN => 
                           n16099);
   U10433 : AOI22_X1 port map( A1 => n17143, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_27_7_port, B1 => 
                           n17145, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_7_port, ZN => 
                           n16093);
   U10432 : AOI22_X1 port map( A1 => n17146, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_23_7_port, B1 => 
                           n17147, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_7_port, ZN => 
                           n16094);
   U10431 : AOI22_X1 port map( A1 => n17148, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_21_7_port, B1 => 
                           n17131, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_7_port, ZN => 
                           n16095);
   U10430 : AOI22_X1 port map( A1 => n17128, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_19_7_port, B1 => 
                           n17134, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_7_port, ZN => 
                           n16096);
   U10429 : NAND4_X1 port map( A1 => n16093, A2 => n16094, A3 => n16095, A4 => 
                           n16096, ZN => n16082);
   U10428 : AOI22_X1 port map( A1 => n17141, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_17_7_port, B1 => 
                           n17341, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_7_port, ZN => 
                           n16089);
   U10427 : AOI22_X1 port map( A1 => n17388, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_9_7_port, B1 => 
                           n17139, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_2_7_port, ZN => 
                           n16090);
   U10426 : AOI22_X1 port map( A1 => n17136, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_12_7_port, B1 => 
                           n17389, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_11_7_port, ZN => 
                           n16091);
   U10425 : AOI22_X1 port map( A1 => n17140, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_14_7_port, B1 => 
                           n17390, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_7_port, ZN => 
                           n16092);
   U10424 : NAND4_X1 port map( A1 => n16089, A2 => n16090, A3 => n16091, A4 => 
                           n16092, ZN => n16083);
   U10423 : AOI22_X1 port map( A1 => n17133, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_7_port, B1 => 
                           n17392, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_4_7_port, ZN => 
                           n16085);
   U10422 : AOI22_X1 port map( A1 => n17334, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_7_port, B1 => 
                           n17144, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_7_port, ZN => 
                           n16086);
   U10421 : AOI22_X1 port map( A1 => n17338, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_6_7_port, B1 => 
                           n17142, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_7_port, ZN => 
                           n16087);
   U10420 : AOI22_X1 port map( A1 => n17336, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_7_port, B1 => 
                           n17391, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_7_port, ZN => 
                           n16088);
   U10419 : NAND4_X1 port map( A1 => n16085, A2 => n16086, A3 => n16087, A4 => 
                           n16088, ZN => n16084);
   U10418 : NOR4_X1 port map( A1 => n16081, A2 => n16082, A3 => n16083, A4 => 
                           n16084, ZN => n14931);
   U10417 : NAND4_X1 port map( A1 => n14925, A2 => n14927, A3 => n14929, A4 => 
                           n14931, ZN => n16003);
   U10416 : AOI22_X1 port map( A1 => n15940, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_31_14_port, B1 => 
                           n15941, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_14_port, ZN => 
                           n16078);
   U10415 : AOI22_X1 port map( A1 => n15938, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_29_14_port, B1 => 
                           n15939, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_14_port, ZN => 
                           n16079);
   U10414 : AOI222_X1 port map( A1 => n15935, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_8_14_port, B1 => 
                           n15936, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_14_port, C1 => 
                           n15937, C2 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_14_port, ZN => 
                           n16080);
   U10413 : AOI22_X1 port map( A1 => n15930, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_27_14_port, B1 => 
                           n15931, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_14_port, ZN => 
                           n16074);
   U10412 : AOI22_X1 port map( A1 => n15928, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_23_14_port, B1 => 
                           n15929, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_14_port, ZN => 
                           n16075);
   U10411 : AOI22_X1 port map( A1 => n15926, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_21_14_port, B1 => 
                           n15927, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_14_port, ZN => 
                           n16076);
   U10410 : AOI22_X1 port map( A1 => n15924, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_19_14_port, B1 => 
                           n15925, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_14_port, ZN => 
                           n16077);
   U10409 : NAND4_X1 port map( A1 => n16074, A2 => n16075, A3 => n16076, A4 => 
                           n16077, ZN => n16063);
   U10408 : AOI22_X1 port map( A1 => n15918, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_17_14_port, B1 => 
                           n17341, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_14_port, ZN => 
                           n16070);
   U10407 : AOI22_X1 port map( A1 => n17388, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_9_14_port, B1 => 
                           n15917, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_2_14_port, ZN => 
                           n16071);
   U10406 : AOI22_X1 port map( A1 => n15914, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_12_14_port, B1 => 
                           n17389, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_11_14_port, ZN => 
                           n16072);
   U10405 : AOI22_X1 port map( A1 => n15912, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_14_14_port, B1 => 
                           n17390, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_14_port, ZN => 
                           n16073);
   U10404 : NAND4_X1 port map( A1 => n16070, A2 => n16071, A3 => n16072, A4 => 
                           n16073, ZN => n16064);
   U10403 : AOI22_X1 port map( A1 => n15906, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_14_port, B1 => 
                           n17392, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_4_14_port, ZN => 
                           n16066);
   U10402 : AOI22_X1 port map( A1 => n17334, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_14_port, B1 => 
                           n15905, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_14_port, ZN => 
                           n16067);
   U10401 : AOI22_X1 port map( A1 => n17338, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_6_14_port, B1 => 
                           n15903, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_14_port, ZN => 
                           n16068);
   U10400 : AOI22_X1 port map( A1 => n17336, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_14_port, B1 => 
                           n17391, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_14_port, ZN => 
                           n16069);
   U10399 : NAND4_X1 port map( A1 => n16066, A2 => n16067, A3 => n16068, A4 => 
                           n16069, ZN => n16065);
   U10398 : NOR4_X1 port map( A1 => n16062, A2 => n16063, A3 => n16064, A4 => 
                           n16065, ZN => n14917);
   U10397 : AOI22_X1 port map( A1 => n17137, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_31_13_port, B1 => 
                           n17138, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_13_port, ZN => 
                           n16059);
   U10396 : AOI22_X1 port map( A1 => n17130, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_29_13_port, B1 => 
                           n17129, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_13_port, ZN => 
                           n16060);
   U10395 : AOI222_X1 port map( A1 => n17135, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_8_13_port, B1 => 
                           n17132, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_13_port, C1 => 
                           n17127, C2 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_13_port, ZN => 
                           n16061);
   U10394 : AOI22_X1 port map( A1 => n17143, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_27_13_port, B1 => 
                           n17145, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_13_port, ZN => 
                           n16055);
   U10393 : AOI22_X1 port map( A1 => n17146, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_23_13_port, B1 => 
                           n17147, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_13_port, ZN => 
                           n16056);
   U10392 : AOI22_X1 port map( A1 => n17148, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_21_13_port, B1 => 
                           n17131, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_13_port, ZN => 
                           n16057);
   U10391 : AOI22_X1 port map( A1 => n17128, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_19_13_port, B1 => 
                           n17134, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_13_port, ZN => 
                           n16058);
   U10390 : NAND4_X1 port map( A1 => n16055, A2 => n16056, A3 => n16057, A4 => 
                           n16058, ZN => n16044);
   U10389 : AOI22_X1 port map( A1 => n17141, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_17_13_port, B1 => 
                           n17341, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_13_port, ZN => 
                           n16051);
   U10388 : AOI22_X1 port map( A1 => n17388, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_9_13_port, B1 => 
                           n17139, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_2_13_port, ZN => 
                           n16052);
   U10387 : AOI22_X1 port map( A1 => n17136, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_12_13_port, B1 => 
                           n17389, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_11_13_port, ZN => 
                           n16053);
   U10386 : AOI22_X1 port map( A1 => n17140, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_14_13_port, B1 => 
                           n17390, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_13_port, ZN => 
                           n16054);
   U10385 : NAND4_X1 port map( A1 => n16051, A2 => n16052, A3 => n16053, A4 => 
                           n16054, ZN => n16045);
   U10384 : AOI22_X1 port map( A1 => n17133, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_13_port, B1 => 
                           n17392, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_4_13_port, ZN => 
                           n16047);
   U10383 : AOI22_X1 port map( A1 => n17334, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_13_port, B1 => 
                           n17144, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_13_port, ZN => 
                           n16048);
   U10382 : AOI22_X1 port map( A1 => n17338, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_6_13_port, B1 => 
                           n17142, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_13_port, ZN => 
                           n16049);
   U10381 : AOI22_X1 port map( A1 => n17336, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_13_port, B1 => 
                           n17391, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_13_port, ZN => 
                           n16050);
   U10380 : NAND4_X1 port map( A1 => n16047, A2 => n16048, A3 => n16049, A4 => 
                           n16050, ZN => n16046);
   U10379 : NOR4_X1 port map( A1 => n16043, A2 => n16044, A3 => n16045, A4 => 
                           n16046, ZN => n14919);
   U10378 : AOI22_X1 port map( A1 => n17137, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_31_12_port, B1 => 
                           n17138, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_12_port, ZN => 
                           n16040);
   U10377 : AOI22_X1 port map( A1 => n17130, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_29_12_port, B1 => 
                           n17129, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_12_port, ZN => 
                           n16041);
   U10376 : AOI222_X1 port map( A1 => n17135, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_8_12_port, B1 => 
                           n17132, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_12_port, C1 => 
                           n17127, C2 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_12_port, ZN => 
                           n16042);
   U10375 : AOI22_X1 port map( A1 => n17143, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_27_12_port, B1 => 
                           n17145, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_12_port, ZN => 
                           n16036);
   U10374 : AOI22_X1 port map( A1 => n17146, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_23_12_port, B1 => 
                           n17147, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_12_port, ZN => 
                           n16037);
   U10373 : AOI22_X1 port map( A1 => n17148, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_21_12_port, B1 => 
                           n17131, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_12_port, ZN => 
                           n16038);
   U10372 : AOI22_X1 port map( A1 => n17128, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_19_12_port, B1 => 
                           n17134, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_12_port, ZN => 
                           n16039);
   U10371 : NAND4_X1 port map( A1 => n16036, A2 => n16037, A3 => n16038, A4 => 
                           n16039, ZN => n16025);
   U10370 : AOI22_X1 port map( A1 => n17141, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_17_12_port, B1 => 
                           n17341, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_12_port, ZN => 
                           n16032);
   U10369 : AOI22_X1 port map( A1 => n17388, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_9_12_port, B1 => 
                           n17139, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_2_12_port, ZN => 
                           n16033);
   U10368 : AOI22_X1 port map( A1 => n17136, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_12_12_port, B1 => 
                           n17389, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_11_12_port, ZN => 
                           n16034);
   U10367 : AOI22_X1 port map( A1 => n17140, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_14_12_port, B1 => 
                           n17390, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_12_port, ZN => 
                           n16035);
   U10366 : NAND4_X1 port map( A1 => n16032, A2 => n16033, A3 => n16034, A4 => 
                           n16035, ZN => n16026);
   U10365 : AOI22_X1 port map( A1 => n17133, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_12_port, B1 => 
                           n17392, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_4_12_port, ZN => 
                           n16028);
   U10364 : AOI22_X1 port map( A1 => n17334, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_12_port, B1 => 
                           n17144, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_12_port, ZN => 
                           n16029);
   U10363 : AOI22_X1 port map( A1 => n17338, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_6_12_port, B1 => 
                           n17142, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_12_port, ZN => 
                           n16030);
   U10362 : AOI22_X1 port map( A1 => n17336, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_12_port, B1 => 
                           n17391, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_12_port, ZN => 
                           n16031);
   U10361 : NAND4_X1 port map( A1 => n16028, A2 => n16029, A3 => n16030, A4 => 
                           n16031, ZN => n16027);
   U10360 : NOR4_X1 port map( A1 => n16024, A2 => n16025, A3 => n16026, A4 => 
                           n16027, ZN => n14921);
   U10359 : AOI22_X1 port map( A1 => n17137, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_31_11_port, B1 => 
                           n17138, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_11_port, ZN => 
                           n16021);
   U10358 : AOI22_X1 port map( A1 => n17130, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_29_11_port, B1 => 
                           n17129, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_11_port, ZN => 
                           n16022);
   U10357 : AOI222_X1 port map( A1 => n17135, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_8_11_port, B1 => 
                           n17132, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_11_port, C1 => 
                           n17127, C2 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_11_port, ZN => 
                           n16023);
   U10356 : AOI22_X1 port map( A1 => n17143, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_27_11_port, B1 => 
                           n17145, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_11_port, ZN => 
                           n16017);
   U10355 : AOI22_X1 port map( A1 => n17146, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_23_11_port, B1 => 
                           n17147, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_11_port, ZN => 
                           n16018);
   U10354 : AOI22_X1 port map( A1 => n17148, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_21_11_port, B1 => 
                           n17131, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_11_port, ZN => 
                           n16019);
   U10353 : AOI22_X1 port map( A1 => n17128, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_19_11_port, B1 => 
                           n17134, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_11_port, ZN => 
                           n16020);
   U10352 : NAND4_X1 port map( A1 => n16017, A2 => n16018, A3 => n16019, A4 => 
                           n16020, ZN => n16006);
   U10351 : AOI22_X1 port map( A1 => n17141, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_17_11_port, B1 => 
                           n17342, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_11_port, ZN => 
                           n16013);
   U10350 : AOI22_X1 port map( A1 => n17388, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_9_11_port, B1 => 
                           n17139, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_2_11_port, ZN => 
                           n16014);
   U10349 : AOI22_X1 port map( A1 => n17136, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_12_11_port, B1 => 
                           n17389, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_11_11_port, ZN => 
                           n16015);
   U10348 : AOI22_X1 port map( A1 => n17140, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_14_11_port, B1 => 
                           n17390, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_11_port, ZN => 
                           n16016);
   U10347 : NAND4_X1 port map( A1 => n16013, A2 => n16014, A3 => n16015, A4 => 
                           n16016, ZN => n16007);
   U10346 : AOI22_X1 port map( A1 => n17133, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_11_port, B1 => 
                           n17392, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_4_11_port, ZN => 
                           n16009);
   U10345 : AOI22_X1 port map( A1 => n17335, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_11_port, B1 => 
                           n17144, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_11_port, ZN => 
                           n16010);
   U10344 : AOI22_X1 port map( A1 => n17339, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_6_11_port, B1 => 
                           n17142, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_11_port, ZN => 
                           n16011);
   U10343 : AOI22_X1 port map( A1 => n17337, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_11_port, B1 => 
                           n17391, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_11_port, ZN => 
                           n16012);
   U10342 : NAND4_X1 port map( A1 => n16009, A2 => n16010, A3 => n16011, A4 => 
                           n16012, ZN => n16008);
   U10341 : NOR4_X1 port map( A1 => n16005, A2 => n16006, A3 => n16007, A4 => 
                           n16008, ZN => n14923);
   U10340 : NAND4_X1 port map( A1 => n14917, A2 => n14919, A3 => n14921, A4 => 
                           n14923, ZN => n16004);
   U10339 : NOR4_X1 port map( A1 => n16001, A2 => n16002, A3 => n16003, A4 => 
                           n16004, ZN => n16000);
   U10338 : NAND4_X1 port map( A1 => n14933, A2 => n14935, A3 => n15999, A4 => 
                           n16000, ZN => n15890);
   U10337 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_31_30_port
                           , A2 => n17137, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_30_port, B2 => 
                           n17138, ZN => n15996);
   U10336 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_29_30_port
                           , A2 => n17130, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_30_port, B2 => 
                           n17129, ZN => n15997);
   U10335 : AOI222_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_8_30_port
                           , A2 => n17135, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_30_port, B2 => 
                           n17132, C1 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_30_port, C2 => 
                           n17127, ZN => n15998);
   U10334 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_27_30_port
                           , A2 => n17143, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_30_port, B2 => 
                           n17145, ZN => n15992);
   U10333 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_23_30_port
                           , A2 => n17146, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_30_port, B2 => 
                           n17147, ZN => n15993);
   U10332 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_21_30_port
                           , A2 => n17148, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_30_port, B2 => 
                           n17131, ZN => n15994);
   U10331 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_19_30_port
                           , A2 => n17128, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_30_port, B2 => 
                           n17134, ZN => n15995);
   U10330 : NAND4_X1 port map( A1 => n15992, A2 => n15993, A3 => n15994, A4 => 
                           n15995, ZN => n15981);
   U10329 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_17_30_port
                           , A2 => n17141, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_30_port, B2 => 
                           n17341, ZN => n15988);
   U10328 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_9_30_port,
                           A2 => n17388, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_2_30_port, B2 => 
                           n17139, ZN => n15989);
   U10327 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_12_30_port
                           , A2 => n17136, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_11_30_port, B2 => 
                           n17389, ZN => n15990);
   U10326 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_14_30_port
                           , A2 => n17140, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_30_port, B2 => 
                           n17390, ZN => n15991);
   U10325 : NAND4_X1 port map( A1 => n15988, A2 => n15989, A3 => n15990, A4 => 
                           n15991, ZN => n15982);
   U10324 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_13_30_port
                           , A2 => n17133, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_4_30_port, B2 => 
                           n17392, ZN => n15984);
   U10323 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_10_30_port
                           , A2 => n17334, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_30_port, B2 => 
                           n17144, ZN => n15985);
   U10322 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_6_30_port,
                           A2 => n17338, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_30_port, B2 => 
                           n17142, ZN => n15986);
   U10321 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_5_30_port,
                           A2 => n17336, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_30_port, B2 => 
                           n17391, ZN => n15987);
   U10320 : NAND4_X1 port map( A1 => n15984, A2 => n15985, A3 => n15986, A4 => 
                           n15987, ZN => n15983);
   U10319 : NOR4_X1 port map( A1 => n15980, A2 => n15981, A3 => n15982, A4 => 
                           n15983, ZN => n14885);
   U10318 : AOI22_X1 port map( A1 => n15940, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_31_29_port, B1 => 
                           n15941, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_29_port, ZN => 
                           n15977);
   U10317 : AOI22_X1 port map( A1 => n15938, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_29_29_port, B1 => 
                           n15939, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_29_port, ZN => 
                           n15978);
   U10316 : AOI222_X1 port map( A1 => n15935, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_8_29_port, B1 => 
                           n15936, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_29_port, C1 => 
                           n15937, C2 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_29_port, ZN => 
                           n15979);
   U10315 : AOI22_X1 port map( A1 => n15930, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_27_29_port, B1 => 
                           n15931, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_29_port, ZN => 
                           n15973);
   U10314 : AOI22_X1 port map( A1 => n15928, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_23_29_port, B1 => 
                           n15929, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_29_port, ZN => 
                           n15974);
   U10313 : AOI22_X1 port map( A1 => n15926, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_21_29_port, B1 => 
                           n15927, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_29_port, ZN => 
                           n15975);
   U10312 : AOI22_X1 port map( A1 => n15924, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_19_29_port, B1 => 
                           n15925, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_29_port, ZN => 
                           n15976);
   U10311 : NAND4_X1 port map( A1 => n15973, A2 => n15974, A3 => n15975, A4 => 
                           n15976, ZN => n15962);
   U10310 : AOI22_X1 port map( A1 => n15918, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_17_29_port, B1 => 
                           n17342, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_29_port, ZN => 
                           n15969);
   U10309 : AOI22_X1 port map( A1 => n17388, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_9_29_port, B1 => 
                           n15917, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_2_29_port, ZN => 
                           n15970);
   U10308 : AOI22_X1 port map( A1 => n15914, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_12_29_port, B1 => 
                           n17389, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_11_29_port, ZN => 
                           n15971);
   U10307 : AOI22_X1 port map( A1 => n15912, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_14_29_port, B1 => 
                           n17390, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_29_port, ZN => 
                           n15972);
   U10306 : NAND4_X1 port map( A1 => n15969, A2 => n15970, A3 => n15971, A4 => 
                           n15972, ZN => n15963);
   U10305 : AOI22_X1 port map( A1 => n15906, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_29_port, B1 => 
                           n17392, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_4_29_port, ZN => 
                           n15965);
   U10304 : AOI22_X1 port map( A1 => n17335, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_29_port, B1 => 
                           n15905, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_29_port, ZN => 
                           n15966);
   U10303 : AOI22_X1 port map( A1 => n17339, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_6_29_port, B1 => 
                           n15903, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_29_port, ZN => 
                           n15967);
   U10302 : AOI22_X1 port map( A1 => n17337, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_29_port, B1 => 
                           n17391, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_29_port, ZN => 
                           n15968);
   U10301 : NAND4_X1 port map( A1 => n15965, A2 => n15966, A3 => n15967, A4 => 
                           n15968, ZN => n15964);
   U10300 : NOR4_X1 port map( A1 => n15961, A2 => n15962, A3 => n15963, A4 => 
                           n15964, ZN => n14887);
   U10299 : AOI22_X1 port map( A1 => n17137, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_31_28_port, B1 => 
                           n17138, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_28_port, ZN => 
                           n15958);
   U10298 : AOI22_X1 port map( A1 => n17130, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_29_28_port, B1 => 
                           n17129, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_28_port, ZN => 
                           n15959);
   U10297 : AOI222_X1 port map( A1 => n17135, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_8_28_port, B1 => 
                           n17132, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_28_port, C1 => 
                           n17127, C2 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_28_port, ZN => 
                           n15960);
   U10296 : AOI22_X1 port map( A1 => n17143, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_27_28_port, B1 => 
                           n17145, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_28_port, ZN => 
                           n15954);
   U10295 : AOI22_X1 port map( A1 => n17146, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_23_28_port, B1 => 
                           n17147, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_28_port, ZN => 
                           n15955);
   U10294 : AOI22_X1 port map( A1 => n17148, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_21_28_port, B1 => 
                           n17131, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_28_port, ZN => 
                           n15956);
   U10293 : AOI22_X1 port map( A1 => n17128, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_19_28_port, B1 => 
                           n17134, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_28_port, ZN => 
                           n15957);
   U10292 : NAND4_X1 port map( A1 => n15954, A2 => n15955, A3 => n15956, A4 => 
                           n15957, ZN => n15943);
   U10291 : AOI22_X1 port map( A1 => n17141, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_17_28_port, B1 => 
                           n17342, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_28_port, ZN => 
                           n15950);
   U10290 : AOI22_X1 port map( A1 => n17388, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_9_28_port, B1 => 
                           n17139, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_2_28_port, ZN => 
                           n15951);
   U10289 : AOI22_X1 port map( A1 => n17136, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_12_28_port, B1 => 
                           n17389, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_11_28_port, ZN => 
                           n15952);
   U10288 : AOI22_X1 port map( A1 => n17140, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_14_28_port, B1 => 
                           n17390, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_28_port, ZN => 
                           n15953);
   U10287 : NAND4_X1 port map( A1 => n15950, A2 => n15951, A3 => n15952, A4 => 
                           n15953, ZN => n15944);
   U10286 : AOI22_X1 port map( A1 => n17133, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_28_port, B1 => 
                           n17392, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_4_28_port, ZN => 
                           n15946);
   U10285 : AOI22_X1 port map( A1 => n17335, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_28_port, B1 => 
                           n17144, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_28_port, ZN => 
                           n15947);
   U10284 : AOI22_X1 port map( A1 => n17339, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_6_28_port, B1 => 
                           n17142, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_28_port, ZN => 
                           n15948);
   U10283 : AOI22_X1 port map( A1 => n17337, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_28_port, B1 => 
                           n17391, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_28_port, ZN => 
                           n15949);
   U10282 : NAND4_X1 port map( A1 => n15946, A2 => n15947, A3 => n15948, A4 => 
                           n15949, ZN => n15945);
   U10281 : NOR4_X1 port map( A1 => n15942, A2 => n15943, A3 => n15944, A4 => 
                           n15945, ZN => n14889);
   U10280 : AOI22_X1 port map( A1 => n17137, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_31_27_port, B1 => 
                           n17138, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_27_port, ZN => 
                           n15932);
   U10279 : AOI22_X1 port map( A1 => n17130, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_29_27_port, B1 => 
                           n17129, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_27_port, ZN => 
                           n15933);
   U10278 : AOI222_X1 port map( A1 => n17135, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_8_27_port, B1 => 
                           n17132, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_27_port, C1 => 
                           n17127, C2 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_27_port, ZN => 
                           n15934);
   U10277 : AOI22_X1 port map( A1 => n17143, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_27_27_port, B1 => 
                           n17145, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_27_port, ZN => 
                           n15920);
   U10276 : AOI22_X1 port map( A1 => n17146, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_23_27_port, B1 => 
                           n17147, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_27_port, ZN => 
                           n15921);
   U10275 : AOI22_X1 port map( A1 => n17148, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_21_27_port, B1 => 
                           n17131, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_27_port, ZN => 
                           n15922);
   U10274 : AOI22_X1 port map( A1 => n17128, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_19_27_port, B1 => 
                           n17134, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_27_port, ZN => 
                           n15923);
   U10273 : NAND4_X1 port map( A1 => n15920, A2 => n15921, A3 => n15922, A4 => 
                           n15923, ZN => n15893);
   U10272 : AOI22_X1 port map( A1 => n17141, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_17_27_port, B1 => 
                           n17342, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_27_port, ZN => 
                           n15908);
   U10271 : AOI22_X1 port map( A1 => n15916, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_9_27_port, B1 => 
                           n17139, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_2_27_port, ZN => 
                           n15909);
   U10270 : AOI22_X1 port map( A1 => n17136, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_12_27_port, B1 => 
                           n15915, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_11_27_port, ZN => 
                           n15910);
   U10269 : AOI22_X1 port map( A1 => n17140, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_14_27_port, B1 => 
                           n15913, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_27_port, ZN => 
                           n15911);
   U10268 : NAND4_X1 port map( A1 => n15908, A2 => n15909, A3 => n15910, A4 => 
                           n15911, ZN => n15894);
   U10267 : AOI22_X1 port map( A1 => n17133, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_27_port, B1 => 
                           n15907, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_4_27_port, ZN => 
                           n15896);
   U10266 : AOI22_X1 port map( A1 => n17335, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_27_port, B1 => 
                           n17144, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_27_port, ZN => 
                           n15897);
   U10265 : AOI22_X1 port map( A1 => n17339, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_6_27_port, B1 => 
                           n17142, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_27_port, ZN => 
                           n15898);
   U10264 : AOI22_X1 port map( A1 => n17337, A2 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_27_port, B1 => 
                           n15901, B2 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_27_port, ZN => 
                           n15899);
   U10263 : NAND4_X1 port map( A1 => n15896, A2 => n15897, A3 => n15898, A4 => 
                           n15899, ZN => n15895);
   U10262 : NOR4_X1 port map( A1 => n15892, A2 => n15893, A3 => n15894, A4 => 
                           n15895, ZN => n14891);
   U10261 : NAND4_X1 port map( A1 => n14885, A2 => n14887, A3 => n14889, A4 => 
                           n14891, ZN => n15891);
   U10259 : NAND4_X1 port map( A1 => n17423, A2 => n17363, A3 => n17322, A4 => 
                           n17310, ZN => n15866);
   U10258 : NAND4_X1 port map( A1 => n17427, A2 => n17324, A3 => n17366, A4 => 
                           n17311, ZN => n15867);
   U10257 : NAND4_X1 port map( A1 => n17344, A2 => n17319, A3 => n17307, A4 => 
                           n17395, ZN => n15868);
   U10256 : NAND4_X1 port map( A1 => n17309, A2 => n17364, A3 => n17323, A4 => 
                           n17426, ZN => n15869);
   U10255 : NOR4_X1 port map( A1 => n15866, A2 => n15867, A3 => n15868, A4 => 
                           n15869, ZN => n15844);
   U10254 : NAND4_X1 port map( A1 => n17394, A2 => n17343, A3 => n17318, A4 => 
                           n17305, ZN => n15846);
   U10253 : NAND4_X1 port map( A1 => n17396, A2 => n17369, A3 => n17321, A4 => 
                           n17306, ZN => n15847);
   U10252 : NAND4_X1 port map( A1 => n17424, A2 => n17325, A3 => n17312, A4 => 
                           n17365, ZN => n15848);
   U10251 : NAND4_X1 port map( A1 => n17425, A2 => n17320, A3 => n17308, A4 => 
                           n17362, ZN => n15849);
   U10250 : NOR4_X1 port map( A1 => n15846, A2 => n15847, A3 => n15848, A4 => 
                           n15849, ZN => n15845);
   U10245 : NAND2_X1 port map( A1 => pipeline_inst_IFID_DEC_26_port, A2 => 
                           n17347, ZN => n14059);
   U10241 : NAND2_X1 port map( A1 => n14126, A2 => n14167, ZN => n15840);
   U10238 : NOR3_X1 port map( A1 => Rst, A2 => n14176, A3 => n14186, ZN => 
                           n14125);
   U11431 : XNOR2_X1 port map( A => pipeline_regDst_to_mem_0_port, B => 
                           pipeline_Reg2_Addr_to_exe_0_port, ZN => n16789);
   U11423 : OAI221_X1 port map( B1 => n17304, B2 => 
                           pipeline_Reg2_Addr_to_exe_1_port, C1 => n17386, C2 
                           => pipeline_Reg2_Addr_to_exe_4_port, A => n16784, ZN
                           => n16779);
   U11321 : NOR2_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_0_port, A2
                           => n13877, ZN => n16731);
   U11320 : AOI22_X1 port map( A1 => n16607, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_13_port, B1 => n17670, 
                           B2 => pipeline_data_to_RF_from_WB_13_port, ZN => 
                           n16732);
   U11319 : OAI21_X1 port map( B1 => n17120, B2 => n16731, A => n16732, ZN => 
                           n16730);
   U11318 : OAI21_X1 port map( B1 => pipeline_immediate_to_exe_13_port, B2 => 
                           n17327, A => n16730, ZN => n15427);
   U11316 : XNOR2_X1 port map( A => n17381, B => n15426, ZN => n16659);
   U11466 : XNOR2_X1 port map( A => n17645, B => 
                           pipeline_Reg1_Addr_to_exe_1_port, ZN => n16808);
   U11465 : NOR2_X1 port map( A1 => n16808, A2 => n16809, ZN => n16807);
   U11472 : XNOR2_X1 port map( A => n17646, B => 
                           pipeline_Reg1_Addr_to_exe_2_port, ZN => n16795);
   U11314 : AOI22_X1 port map( A1 => n17663, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_13_port, B1 => n17664, 
                           B2 => n13958, ZN => n16729);
   U11312 : NAND2_X1 port map( A1 => n16659, A2 => 
                           pipeline_stageE_input1_to_ALU_13_port, ZN => n15416)
                           ;
   U11233 : NAND2_X1 port map( A1 => n16691, A2 => n12649, ZN => n15053);
   U11230 : AOI22_X1 port map( A1 => n17663, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_3_port, B1 => n17664, 
                           B2 => n13844, ZN => n16689);
   U11227 : NOR2_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_0_port, A2
                           => n13838, ZN => n16685);
   U11226 : AOI22_X1 port map( A1 => n16607, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_4_port, B1 => n15123, 
                           B2 => pipeline_data_to_RF_from_WB_4_port, ZN => 
                           n16686);
   U11225 : NOR2_X1 port map( A1 => pipeline_immediate_to_exe_4_port, A2 => 
                           n17327, ZN => n16687);
   U11224 : AOI221_X1 port map( B1 => n16685, B2 => n16686, C1 => n17120, C2 =>
                           n16686, A => n16687, ZN => n4376);
   U11222 : OAI22_X1 port map( A1 => n17381, A2 => n17737, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, B2 
                           => pipeline_stageE_EXE_ALU_add_alu_sCout_0_port, ZN 
                           => n16683);
   U11220 : AOI22_X1 port map( A1 => n17663, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_4_port, B1 => n17664, 
                           B2 => n13836, ZN => n16684);
   U11215 : NAND2_X1 port map( A1 => n15564, A2 => n16683, ZN => n15568);
   U11279 : NOR2_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_0_port, A2
                           => n13834, ZN => n16711);
   U11278 : AOI22_X1 port map( A1 => n16607, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_5_port, B1 => n17670, 
                           B2 => pipeline_data_to_RF_from_WB_5_port, ZN => 
                           n16712);
   U11277 : OAI21_X1 port map( B1 => n17120, B2 => n16711, A => n16712, ZN => 
                           n16710);
   U11276 : OAI21_X1 port map( B1 => pipeline_immediate_to_exe_5_port, B2 => 
                           n17327, A => n16710, ZN => n15553);
   U11272 : NOR2_X1 port map( A1 => n16677, A2 => 
                           pipeline_stageE_input1_to_ALU_5_port, ZN => n15542);
   U11213 : NOR2_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_0_port, A2
                           => n13843, ZN => n16680);
   U11212 : AOI22_X1 port map( A1 => n17665, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_6_port, B1 => n17123, 
                           B2 => pipeline_data_to_RF_from_WB_6_port, ZN => 
                           n16681);
   U11211 : OAI21_X1 port map( B1 => n17120, B2 => n16680, A => n16681, ZN => 
                           n16679);
   U11210 : OAI21_X1 port map( B1 => pipeline_immediate_to_exe_6_port, B2 => 
                           n17327, A => n16679, ZN => n15538);
   U11208 : XNOR2_X1 port map( A => n17381, B => n15537, ZN => n16676);
   U11206 : AOI22_X1 port map( A1 => n17663, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_6_port, B1 => n17664, 
                           B2 => n13842, ZN => n16678);
   U11204 : NAND2_X1 port map( A1 => n16676, A2 => 
                           pipeline_stageE_input1_to_ALU_6_port, ZN => n15525);
   U11203 : NAND2_X1 port map( A1 => n16677, A2 => 
                           pipeline_stageE_input1_to_ALU_5_port, ZN => n15540);
   U11281 : AOI22_X1 port map( A1 => n17663, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_7_port, B1 => n17664, 
                           B2 => n13839, ZN => n16713);
   U11286 : NOR2_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_0_port, A2
                           => n13841, ZN => n16715);
   U11285 : AOI22_X1 port map( A1 => n16607, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_7_port, B1 => n17670, 
                           B2 => pipeline_data_to_RF_from_WB_7_port, ZN => 
                           n16716);
   U11284 : OAI21_X1 port map( B1 => n17120, B2 => n16715, A => n16716, ZN => 
                           n16714);
   U11283 : OAI21_X1 port map( B1 => pipeline_immediate_to_exe_7_port, B2 => 
                           n17327, A => n16714, ZN => n15512);
   U11293 : NOR2_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_0_port, A2
                           => n13875, ZN => n16718);
   U11292 : AOI22_X1 port map( A1 => n16607, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_8_port, B1 => n17670, 
                           B2 => pipeline_data_to_RF_from_WB_8_port, ZN => 
                           n16719);
   U11291 : OAI21_X1 port map( B1 => n17120, B2 => n16718, A => n16719, ZN => 
                           n16717);
   U11290 : OAI21_X1 port map( B1 => pipeline_immediate_to_exe_8_port, B2 => 
                           n17327, A => n16717, ZN => n15498);
   U11288 : XNOR2_X1 port map( A => n17381, B => n15505, ZN => n16672);
   U11196 : NAND2_X1 port map( A1 => n16672, A2 => 
                           pipeline_stageE_input1_to_ALU_8_port, ZN => n15479);
   U11191 : NOR2_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_0_port, A2
                           => n13822, ZN => n16669);
   U11190 : AOI22_X1 port map( A1 => n17665, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_9_port, B1 => n17123, 
                           B2 => pipeline_data_to_RF_from_WB_9_port, ZN => 
                           n16670);
   U11189 : OAI21_X1 port map( B1 => n17120, B2 => n16669, A => n16670, ZN => 
                           n16668);
   U11188 : OAI21_X1 port map( B1 => pipeline_immediate_to_exe_9_port, B2 => 
                           n17327, A => n16668, ZN => n15492);
   U11186 : XNOR2_X1 port map( A => n17381, B => n15491, ZN => n16667);
   U11185 : NOR2_X1 port map( A1 => pipeline_stageE_input1_to_ALU_9_port, A2 =>
                           n16667, ZN => n15477);
   U11304 : NOR2_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_0_port, A2
                           => n13827, ZN => n16723);
   U11303 : AOI22_X1 port map( A1 => n17665, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_10_port, B1 => n17670, 
                           B2 => pipeline_data_to_RF_from_WB_10_port, ZN => 
                           n16724);
   U11302 : OAI21_X1 port map( B1 => n17120, B2 => n16723, A => n16724, ZN => 
                           n16722);
   U11301 : OAI21_X1 port map( B1 => pipeline_immediate_to_exe_10_port, B2 => 
                           n17327, A => n16722, ZN => n15474);
   U11299 : AOI22_X1 port map( A1 => n17663, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_10_port, B1 => n17664, 
                           B2 => n13826, ZN => n16721);
   U11181 : NAND2_X1 port map( A1 => n16666, A2 => 
                           pipeline_stageE_input1_to_ALU_10_port, ZN => n15463)
                           ;
   U11182 : NAND2_X1 port map( A1 => n16667, A2 => 
                           pipeline_stageE_input1_to_ALU_9_port, ZN => n15480);
   U11306 : AOI22_X1 port map( A1 => n17663, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_11_port, B1 => n17664, 
                           B2 => n13823, ZN => n16725);
   U11311 : NOR2_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_0_port, A2
                           => n13825, ZN => n16727);
   U11310 : AOI22_X1 port map( A1 => n16607, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_11_port, B1 => n17670, 
                           B2 => pipeline_data_to_RF_from_WB_11_port, ZN => 
                           n16728);
   U11309 : OAI21_X1 port map( B1 => n17120, B2 => n16727, A => n16728, ZN => 
                           n16726);
   U11308 : OAI21_X1 port map( B1 => pipeline_immediate_to_exe_11_port, B2 => 
                           n17327, A => n16726, ZN => n15449);
   U11178 : NOR2_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_0_port, A2
                           => n13815, ZN => n16662);
   U11176 : OAI21_X1 port map( B1 => n17120, B2 => n16662, A => n16663, ZN => 
                           n16661);
   U11175 : OAI21_X1 port map( B1 => pipeline_immediate_to_exe_12_port, B2 => 
                           n17327, A => n16661, ZN => n15435);
   U11173 : XNOR2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_add_alu_sCout_0_port, B => 
                           n15442, ZN => n16658);
   U11171 : AOI22_X1 port map( A1 => n17663, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_12_port, B1 => n17664, 
                           B2 => n13814, ZN => n16660);
   U11168 : NOR2_X1 port map( A1 => n16658, A2 => n17080, ZN => n15431);
   U11165 : NOR2_X1 port map( A1 => pipeline_stageE_input1_to_ALU_13_port, A2 
                           => n16659, ZN => n15414);
   U11163 : NAND2_X1 port map( A1 => n17080, A2 => n16658, ZN => n15430);
   U11162 : NOR2_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_0_port, A2
                           => n13874, ZN => n16655);
   U11161 : AOI22_X1 port map( A1 => n17665, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_14_port, B1 => n17670, 
                           B2 => pipeline_data_to_RF_from_WB_14_port, ZN => 
                           n16656);
   U11160 : OAI21_X1 port map( B1 => n17120, B2 => n16655, A => n16656, ZN => 
                           n16654);
   U11159 : OAI21_X1 port map( B1 => pipeline_immediate_to_exe_14_port, B2 => 
                           n17327, A => n16654, ZN => n15411);
   U11157 : XNOR2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_add_alu_sCout_0_port, B => 
                           n15410, ZN => n16651);
   U11155 : AOI22_X1 port map( A1 => n17663, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_14_port, B1 => n17664, 
                           B2 => n13960, ZN => n16653);
   U11152 : NAND2_X1 port map( A1 => n16651, A2 => n17100, ZN => n15400);
   U11149 : NOR2_X1 port map( A1 => n17100, A2 => n16651, ZN => n15398);
   U11147 : NOR2_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_0_port, A2
                           => n13878, ZN => n16648);
   U11146 : AOI22_X1 port map( A1 => n17665, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_15_port, B1 => n17670, 
                           B2 => pipeline_data_to_RF_from_WB_15_port, ZN => 
                           n16649);
   U11145 : OAI21_X1 port map( B1 => n17120, B2 => n16648, A => n16649, ZN => 
                           n16647);
   U11144 : OAI21_X1 port map( B1 => pipeline_immediate_to_exe_15_port, B2 => 
                           n17327, A => n16647, ZN => n15386);
   U11143 : XNOR2_X1 port map( A => n17381, B => n15386, ZN => n15397);
   U11140 : AOI22_X1 port map( A1 => n17663, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_17_port, B1 => n17664, 
                           B2 => n13946, ZN => n16645);
   U11138 : NOR2_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_0_port, A2
                           => n13879, ZN => n16643);
   U11137 : AOI22_X1 port map( A1 => n17665, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_17_port, B1 => n17123, 
                           B2 => pipeline_data_to_RF_from_WB_17_port, ZN => 
                           n16644);
   U11136 : OAI21_X1 port map( B1 => n17120, B2 => n16643, A => n16644, ZN => 
                           n16642);
   U11135 : OAI21_X1 port map( B1 => pipeline_immediate_to_exe_17_port, B2 => 
                           n17327, A => n16642, ZN => n15363);
   U11133 : XNOR2_X1 port map( A => n17381, B => n15362, ZN => n16633);
   U11132 : NOR2_X1 port map( A1 => pipeline_stageE_input1_to_ALU_17_port, A2 
                           => n16633, ZN => n16632);
   U11128 : OAI21_X1 port map( B1 => n17105, B2 => n17426, A => n16641, ZN => 
                           pipeline_stageE_input1_to_ALU_16_port);
   U11127 : NOR2_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_0_port, A2
                           => n13873, ZN => n16639);
   U11125 : OAI21_X1 port map( B1 => n17120, B2 => n16639, A => n16640, ZN => 
                           n16638);
   U11124 : OAI21_X1 port map( B1 => pipeline_immediate_to_exe_16_port, B2 => 
                           n17327, A => n16638, ZN => n15372);
   U11122 : XNOR2_X1 port map( A => n17381, B => n15379, ZN => n15369);
   U11333 : NOR2_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_0_port, A2
                           => n13872, ZN => n16736);
   U11332 : AOI22_X1 port map( A1 => n16607, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_18_port, B1 => n17670, 
                           B2 => pipeline_data_to_RF_from_WB_18_port, ZN => 
                           n16737);
   U11331 : OAI21_X1 port map( B1 => n17120, B2 => n16736, A => n16737, ZN => 
                           n16735);
   U11330 : OAI21_X1 port map( B1 => pipeline_immediate_to_exe_18_port, B2 => 
                           n17327, A => n16735, ZN => n15346);
   U11115 : NOR2_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_0_port, A2
                           => n13880, ZN => n16635);
   U11114 : AOI22_X1 port map( A1 => n17666, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_19_port, B1 => n17670, 
                           B2 => pipeline_data_to_RF_from_WB_19_port, ZN => 
                           n16636);
   U11113 : OAI21_X1 port map( B1 => n17120, B2 => n16635, A => n16636, ZN => 
                           n16634);
   U11112 : OAI21_X1 port map( B1 => pipeline_immediate_to_exe_19_port, B2 => 
                           n17327, A => n16634, ZN => n15331);
   U11110 : XNOR2_X1 port map( A => n17381, B => n15330, ZN => n15314);
   U11100 : NAND2_X1 port map( A1 => n17097, A2 => n15332, ZN => n15316);
   U11349 : NOR2_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_0_port, A2
                           => n13881, ZN => n16744);
   U11348 : AOI22_X1 port map( A1 => n17666, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_21_port, B1 => n17670, 
                           B2 => pipeline_data_to_RF_from_WB_21_port, ZN => 
                           n16745);
   U11347 : OAI21_X1 port map( B1 => n17120, B2 => n16744, A => n16745, ZN => 
                           n16743);
   U11346 : OAI21_X1 port map( B1 => pipeline_immediate_to_exe_21_port, B2 => 
                           n17327, A => n16743, ZN => n15285);
   U11344 : AOI22_X1 port map( A1 => n17663, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_21_port, B1 => n17664, 
                           B2 => n13950, ZN => n16742);
   U11342 : NOR2_X1 port map( A1 => n16626, A2 => 
                           pipeline_stageE_input1_to_ALU_21_port, ZN => n15301)
                           ;
   U11341 : NOR2_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_0_port, A2
                           => n13871, ZN => n16740);
   U11340 : AOI22_X1 port map( A1 => n17666, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_20_port, B1 => n17670, 
                           B2 => pipeline_data_to_RF_from_WB_20_port, ZN => 
                           n16741);
   U11339 : OAI21_X1 port map( B1 => n17120, B2 => n16740, A => n16741, ZN => 
                           n16739);
   U11338 : OAI21_X1 port map( B1 => pipeline_immediate_to_exe_20_port, B2 => 
                           n17327, A => n16739, ZN => n15312);
   U11336 : AOI22_X1 port map( A1 => n17663, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_20_port, B1 => n17664, 
                           B2 => n13949, ZN => n16738);
   U11102 : NOR2_X1 port map( A1 => n16629, A2 => 
                           pipeline_stageE_input1_to_ALU_20_port, ZN => n15298)
                           ;
   U11108 : NAND2_X1 port map( A1 => n15369, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_A_16_port, ZN 
                           => n15382);
   U11107 : NAND2_X1 port map( A1 => n16633, A2 => 
                           pipeline_stageE_input1_to_ALU_17_port, ZN => n15366)
                           ;
   U11106 : OAI21_X1 port map( B1 => n16632, B2 => n15382, A => n15366, ZN => 
                           n15352);
   U11104 : OAI221_X1 port map( B1 => n15352, B2 => n15348, C1 => n15352, C2 =>
                           pipeline_stageE_input1_to_ALU_18_port, A => n16630, 
                           ZN => n15319);
   U11334 : NAND2_X1 port map( A1 => n16629, A2 => 
                           pipeline_stageE_input1_to_ALU_20_port, ZN => n15297)
                           ;
   U11098 : NAND2_X1 port map( A1 => n16626, A2 => 
                           pipeline_stageE_input1_to_ALU_21_port, ZN => n15299)
                           ;
   U11359 : AOI22_X1 port map( A1 => n17663, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_22_port, B1 => n17664, 
                           B2 => n13951, ZN => n16749);
   U11357 : NOR2_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_0_port, A2
                           => n13870, ZN => n16747);
   U11356 : AOI22_X1 port map( A1 => n17666, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_22_port, B1 => n17670, 
                           B2 => pipeline_data_to_RF_from_WB_22_port, ZN => 
                           n16748);
   U11355 : OAI21_X1 port map( B1 => n17120, B2 => n16747, A => n16748, ZN => 
                           n16746);
   U11354 : OAI21_X1 port map( B1 => pipeline_immediate_to_exe_22_port, B2 => 
                           n17327, A => n16746, ZN => n15279);
   U11352 : XNOR2_X1 port map( A => n17381, B => n15278, ZN => n16624);
   U11351 : NAND2_X1 port map( A1 => pipeline_stageE_input1_to_ALU_22_port, A2 
                           => n16624, ZN => n15268);
   U11364 : NOR2_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_0_port, A2
                           => n13882, ZN => n16751);
   U11362 : OAI21_X1 port map( B1 => n17120, B2 => n16751, A => n16752, ZN => 
                           n16750);
   U11361 : OAI21_X1 port map( B1 => pipeline_immediate_to_exe_23_port, B2 => 
                           n17327, A => n16750, ZN => n15261);
   U11095 : NOR2_X1 port map( A1 => n16624, A2 => 
                           pipeline_stageE_input1_to_ALU_22_port, ZN => n15265)
                           ;
   U11090 : AOI22_X1 port map( A1 => n17663, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_24_port, B1 => n17664, 
                           B2 => n13963, ZN => n16618);
   U11087 : NOR2_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_0_port, A2
                           => n13869, ZN => n16615);
   U11086 : AOI22_X1 port map( A1 => n17666, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_24_port, B1 => n17670, 
                           B2 => pipeline_data_to_RF_from_WB_24_port, ZN => 
                           n16616);
   U11085 : OAI21_X1 port map( B1 => n17120, B2 => n16615, A => n16616, ZN => 
                           n16614);
   U11084 : OAI21_X1 port map( B1 => pipeline_immediate_to_exe_24_port, B2 => 
                           n17327, A => n16614, ZN => n15246);
   U11082 : XNOR2_X1 port map( A => n17381, B => n15245, ZN => n15249);
   U11080 : NAND2_X1 port map( A1 => n15249, A2 => 
                           pipeline_stageE_input1_to_ALU_24_port, ZN => n15250)
                           ;
   U11369 : AOI22_X1 port map( A1 => n17663, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_25_port, B1 => n17664, 
                           B2 => n13953, ZN => n16754);
   U11374 : NOR2_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_0_port, A2
                           => n13883, ZN => n16756);
   U11372 : OAI21_X1 port map( B1 => n17120, B2 => n16756, A => n16757, ZN => 
                           n16755);
   U11371 : OAI21_X1 port map( B1 => pipeline_immediate_to_exe_25_port, B2 => 
                           n17327, A => n16755, ZN => n15224);
   U11382 : NOR2_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_0_port, A2
                           => n13868, ZN => n16760);
   U11381 : AOI22_X1 port map( A1 => n17666, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_26_port, B1 => n17123, 
                           B2 => pipeline_data_to_RF_from_WB_26_port, ZN => 
                           n16761);
   U11380 : OAI21_X1 port map( B1 => n17120, B2 => n16760, A => n16761, ZN => 
                           n16759);
   U11379 : OAI21_X1 port map( B1 => pipeline_immediate_to_exe_26_port, B2 => 
                           n17327, A => n16759, ZN => n15216);
   U11377 : AOI22_X1 port map( A1 => n17663, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_26_port, B1 => n17664, 
                           B2 => n13954, ZN => n16758);
   U11375 : NOR2_X1 port map( A1 => n16612, A2 => 
                           pipeline_stageE_input1_to_ALU_26_port, ZN => n15220)
                           ;
   U11077 : NAND2_X1 port map( A1 => n16612, A2 => 
                           pipeline_stageE_input1_to_ALU_26_port, ZN => n15221)
                           ;
   U11384 : AOI22_X1 port map( A1 => n17663, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_27_port, B1 => n17664, 
                           B2 => n13955, ZN => n16762);
   U11389 : NOR2_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_0_port, A2
                           => n13884, ZN => n16764);
   U11388 : AOI22_X1 port map( A1 => n17665, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_27_port, B1 => n17670, 
                           B2 => pipeline_data_to_RF_from_WB_27_port, ZN => 
                           n16765);
   U11387 : OAI21_X1 port map( B1 => n17120, B2 => n16764, A => n16765, ZN => 
                           n16763);
   U11386 : OAI21_X1 port map( B1 => pipeline_immediate_to_exe_27_port, B2 => 
                           n17327, A => n16763, ZN => n15202);
   U11397 : NOR2_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_0_port, A2
                           => n13867, ZN => n16768);
   U11396 : AOI22_X1 port map( A1 => n17665, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_28_port, B1 => n17670, 
                           B2 => pipeline_data_to_RF_from_WB_28_port, ZN => 
                           n16769);
   U11395 : OAI21_X1 port map( B1 => n17120, B2 => n16768, A => n16769, ZN => 
                           n16767);
   U11394 : OAI21_X1 port map( B1 => pipeline_immediate_to_exe_28_port, B2 => 
                           n17327, A => n16767, ZN => n15182);
   U11074 : NAND2_X1 port map( A1 => pipeline_stageE_input1_to_ALU_28_port, A2 
                           => n16611, ZN => n15163);
   U9633 : NAND2_X1 port map( A1 => n15166, A2 => n15163, ZN => n15191);
   U9670 : OAI21_X1 port map( B1 => n15249, B2 => n17158, A => n15250, ZN => 
                           n15247);
   U9652 : NOR2_X1 port map( A1 => n15219, A2 => n15220, ZN => n15217);
   U9680 : OAI21_X1 port map( B1 => n15265, B2 => n15267, A => n15268, ZN => 
                           n15264);
   U9679 : NAND2_X1 port map( A1 => n17092, A2 => n15264, ZN => n15266);
   U9678 : OAI22_X1 port map( A1 => n17092, A2 => n15264, B1 => n15265, B2 => 
                           n15266, ZN => n15262);
   U9724 : NAND2_X1 port map( A1 => n15319, A2 => n15335, ZN => n15334);
   U9691 : NOR2_X1 port map( A1 => n15281, A2 => n15265, ZN => n15280);
   U9690 : XNOR2_X1 port map( A => n15267, B => n15280, ZN => n15024);
   U9661 : XNOR2_X1 port map( A => n15233, B => n17115, ZN => n15020);
   U9702 : NAND2_X1 port map( A1 => n15299, A2 => n15300, ZN => n15294);
   U9715 : NOR2_X1 port map( A1 => n15314, A2 => 
                           pipeline_stageE_input1_to_ALU_19_port, ZN => n15318)
                           ;
   U9714 : NOR2_X1 port map( A1 => n15318, A2 => n15319, ZN => n15317);
   U9701 : AOI21_X1 port map( B1 => n15296, B2 => n15297, A => n15298, ZN => 
                           n15295);
   U9753 : NAND2_X1 port map( A1 => n15382, A2 => n15383, ZN => n15381);
   U9777 : AOI21_X1 port map( B1 => n15429, B2 => n15430, A => n15431, ZN => 
                           n15415);
   U9769 : OAI21_X1 port map( B1 => n15414, B2 => n15415, A => n15416, ZN => 
                           n15399);
   U9761 : OAI21_X1 port map( B1 => n15398, B2 => n15399, A => n15400, ZN => 
                           n15395);
   U9778 : NAND2_X1 port map( A1 => n15432, A2 => n15416, ZN => n15428);
   U9808 : NAND2_X1 port map( A1 => n15463, A2 => n17587, ZN => n15475);
   U9796 : OAI21_X1 port map( B1 => n15461, B2 => n15462, A => n15463, ZN => 
                           n15460);
   U9795 : XNOR2_X1 port map( A => n15459, B => n15460, ZN => n15458);
   U9794 : XNOR2_X1 port map( A => n17082, B => n15458, ZN => n15040);
   U9826 : NAND2_X1 port map( A1 => n15479, A2 => n15509, ZN => n15507);
   U9837 : NAND2_X1 port map( A1 => n15526, A2 => n15527, ZN => n15524);
   U9836 : NAND2_X1 port map( A1 => n15524, A2 => n15525, ZN => n15523);
   U9835 : XNOR2_X1 port map( A => n17089, B => n15523, ZN => n15522);
   U9834 : XNOR2_X1 port map( A => n15521, B => n15522, ZN => n15037);
   U9847 : NAND2_X1 port map( A1 => n15527, A2 => n15525, ZN => n15539);
   U9846 : XNOR2_X1 port map( A => n15526, B => n15539, ZN => n15043);
   U9858 : NOR2_X1 port map( A1 => n15555, A2 => n15542, ZN => n15554);
   U9866 : NAND2_X1 port map( A1 => n15568, A2 => n15569, ZN => n15567);
   U9899 : AOI21_X1 port map( B1 => n15058, B2 => n15053, A => n15055, ZN => 
                           n15592);
   U9896 : AOI21_X1 port map( B1 => n15594, B2 => n15053, A => n15055, ZN => 
                           n15593);
   U9513 : NAND2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_add_alu_sCout_0_port, A2 => 
                           n15058, ZN => n15057);
   U9512 : OAI21_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_add_alu_sCout_0_port, B2 => 
                           n15056, A => n15057, ZN => n15051);
   U9510 : NAND2_X1 port map( A1 => n15053, A2 => n15054, ZN => n15052);
   U9509 : XNOR2_X1 port map( A => n15051, B => n15052, ZN => n14948);
   U9818 : NAND2_X1 port map( A1 => n15480, A2 => n15495, ZN => n15493);
   U9786 : NAND2_X1 port map( A1 => n15430, A2 => n15446, ZN => n15444);
   U9768 : NOR2_X1 port map( A1 => n15413, A2 => n15398, ZN => n15412);
   U9716 : NOR2_X1 port map( A1 => n15320, A2 => n15298, ZN => n15313);
   U9712 : XNOR2_X1 port map( A => n15313, B => n15296, ZN => n15026);
   U11407 : NOR2_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_0_port, A2
                           => n13885, ZN => n16772);
   U11405 : OAI21_X1 port map( B1 => n17120, B2 => n16772, A => n16773, ZN => 
                           n16771);
   U11404 : OAI21_X1 port map( B1 => pipeline_immediate_to_exe_29_port, B2 => 
                           n17327, A => n16771, ZN => n15169);
   U11402 : XNOR2_X1 port map( A => n17381, B => n15176, ZN => n16609);
   U9613 : NAND2_X1 port map( A1 => n15165, A2 => n15166, ZN => n15146);
   U11071 : NAND2_X1 port map( A1 => pipeline_stageE_input1_to_ALU_29_port, A2 
                           => n16609, ZN => n15147);
   U9612 : OAI21_X1 port map( B1 => n15163, B2 => n15164, A => n15147, ZN => 
                           n15162);
   U11415 : NOR2_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_0_port, A2
                           => n13866, ZN => n16775);
   U11414 : AOI22_X1 port map( A1 => n17665, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_30_port, B1 => n17123, 
                           B2 => pipeline_data_to_RF_from_WB_30_port, ZN => 
                           n16776);
   U11413 : OAI21_X1 port map( B1 => n17642, B2 => n16775, A => n16776, ZN => 
                           n16774);
   U11412 : OAI21_X1 port map( B1 => pipeline_immediate_to_exe_30_port, B2 => 
                           n17327, A => n16774, ZN => n15150);
   U11410 : XNOR2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_add_alu_sCout_0_port, B => 
                           n15157, ZN => n16608);
   U11435 : AOI22_X1 port map( A1 => n16619, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_30_port, B1 => n17664, 
                           B2 => n13957, ZN => n16792);
   U11409 : NAND2_X1 port map( A1 => n17083, A2 => n16608, ZN => n15142);
   U9608 : NAND2_X1 port map( A1 => n15138, A2 => n15142, ZN => n15160);
   U11439 : AOI22_X1 port map( A1 => n17663, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_31_port, B1 => n17664, 
                           B2 => n13966, ZN => n16793);
   U11067 : NOR2_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_0_port, A2
                           => n13886, ZN => n16605);
   U11066 : AOI22_X1 port map( A1 => n17666, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_31_port, B1 => n17670, 
                           B2 => pipeline_data_to_RF_from_WB_31_port, ZN => 
                           n16606);
   U11065 : OAI21_X1 port map( B1 => n17642, B2 => n16605, A => n16606, ZN => 
                           n16603);
   U11064 : OAI21_X1 port map( B1 => pipeline_immediate_to_exe_31_port, B2 => 
                           n17327, A => n16603, ZN => n15134);
   U9882 : NOR2_X1 port map( A1 => n17381, A2 => n15586, ZN => n15583);
   U9879 : NAND2_X1 port map( A1 => n15583, A2 => n17405, ZN => n15584);
   U9881 : NAND2_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_3_port, A2
                           => n15583, ZN => n15581);
   U9876 : NAND2_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_2_port, A2
                           => n15583, ZN => n15582);
   U10219 : NOR2_X1 port map( A1 => n15834, A2 => n14127, ZN => n15607);
   U10053 : AOI22_X1 port map( A1 => pipeline_stageF_PC_plus4_N35, A2 => n17108
                           , B1 => n17674, B2 => n13865, ZN => n15689);
   U10051 : AOI22_X1 port map( A1 => pipeline_stageD_target_Jump_temp_28_port, 
                           A2 => n15607, B1 => n17106, B2 => n15692, ZN => 
                           n15690);
   U10050 : AOI22_X1 port map( A1 => pipeline_data_to_RF_from_WB_28_port, A2 =>
                           n17332, B1 => pipeline_Alu_Out_Addr_to_mem_28_port, 
                           B2 => n17330, ZN => n15691);
   U10059 : AOI22_X1 port map( A1 => pipeline_stageF_PC_plus4_N34, A2 => n17108
                           , B1 => n15611, B2 => n13864, ZN => n15694);
   U10057 : AOI22_X1 port map( A1 => pipeline_stageD_target_Jump_temp_27_port, 
                           A2 => n17676, B1 => n17106, B2 => n15697, ZN => 
                           n15695);
   U10056 : AOI22_X1 port map( A1 => pipeline_data_to_RF_from_WB_27_port, A2 =>
                           n17332, B1 => pipeline_Alu_Out_Addr_to_mem_27_port, 
                           B2 => n17330, ZN => n15696);
   U9892 : NAND2_X1 port map( A1 => n17421, A2 => n14995, ZN => n15588);
   U9596 : AOI22_X1 port map( A1 => n17150, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N38, B1 => n17149,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_N70, ZN => 
                           n15128);
   U9595 : AOI22_X1 port map( A1 => n17680, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N168, B1 => n17126
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N136, ZN 
                           => n15129);
   U9594 : AOI22_X1 port map( A1 => n17419, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N233, B1 => n17360
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N265, ZN 
                           => n15130);
   U9593 : NAND4_X1 port map( A1 => n15128, A2 => n15129, A3 => n15130, A4 => 
                           n15131, ZN => n15127);
   U9591 : NAND2_X1 port map( A1 => n15124, A2 => n15125, ZN => 
                           pipeline_EXMEM_stage_N38);
   U9607 : NOR2_X1 port map( A1 => pipeline_stageE_input1_to_ALU_30_port, A2 =>
                           n15150, ZN => n15151);
   U9606 : AOI22_X1 port map( A1 => n17150, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N37, B1 => n17149,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_N69, ZN => 
                           n15154);
   U9605 : AOI22_X1 port map( A1 => n17359, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N167, B1 => n14964
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N135, ZN 
                           => n15155);
   U9604 : AOI22_X1 port map( A1 => n17419, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N232, B1 => n17360
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N264, ZN 
                           => n15156);
   U9603 : AOI211_X1 port map( C1 => n14954, C2 => n15151, A => n15152, B => 
                           n15153, ZN => n15148);
   U9602 : OAI211_X1 port map( C1 => n15009, C2 => n14949, A => n15148, B => 
                           n15149, ZN => pipeline_EXMEM_stage_N37);
   U10065 : AOI22_X1 port map( A1 => pipeline_stageF_PC_plus4_N33, A2 => n17108
                           , B1 => n17674, B2 => n13863, ZN => n15699);
   U10063 : AOI22_X1 port map( A1 => pipeline_stageD_target_Jump_temp_26_port, 
                           A2 => n17676, B1 => n17106, B2 => n15702, ZN => 
                           n15700);
   U10062 : AOI22_X1 port map( A1 => pipeline_data_to_RF_from_WB_26_port, A2 =>
                           n17332, B1 => pipeline_Alu_Out_Addr_to_mem_26_port, 
                           B2 => n17330, ZN => n15701);
   U9620 : NOR2_X1 port map( A1 => pipeline_stageE_input1_to_ALU_29_port, A2 =>
                           n15169, ZN => n15170);
   U9887 : NAND2_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_4_port, A2
                           => n15573, ZN => n14967);
   U9618 : AOI22_X1 port map( A1 => n17150, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N36, B1 => n17149,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_N68, ZN => 
                           n15173);
   U9617 : AOI22_X1 port map( A1 => n17359, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N166, B1 => n17126
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N134, ZN 
                           => n15174);
   U9616 : AOI22_X1 port map( A1 => n17419, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N231, B1 => n17681
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N263, ZN 
                           => n15175);
   U9615 : AOI211_X1 port map( C1 => n14954, C2 => n15170, A => n15171, B => 
                           n15172, ZN => n15167);
   U9614 : OAI211_X1 port map( C1 => n15010, C2 => n14949, A => n15167, B => 
                           n15168, ZN => pipeline_EXMEM_stage_N36);
   U9631 : NOR2_X1 port map( A1 => pipeline_stageE_input1_to_ALU_28_port, A2 =>
                           n15182, ZN => n15183);
   U9628 : AOI22_X1 port map( A1 => n17150, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N35, B1 => n17149,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_N67, ZN => 
                           n15186);
   U9627 : AOI22_X1 port map( A1 => n17359, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N165, B1 => n17126
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N133, ZN 
                           => n15187);
   U9626 : AOI22_X1 port map( A1 => n17419, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N230, B1 => n17681
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N262, ZN 
                           => n15188);
   U9625 : AOI211_X1 port map( C1 => n14954, C2 => n15183, A => n15184, B => 
                           n15185, ZN => n15180);
   U9624 : OAI211_X1 port map( C1 => n15011, C2 => n14949, A => n15180, B => 
                           n15181, ZN => pipeline_EXMEM_stage_N35);
   U10071 : AOI22_X1 port map( A1 => pipeline_stageF_PC_plus4_N32, A2 => n17108
                           , B1 => n17674, B2 => n13862, ZN => n15704);
   U10069 : AOI22_X1 port map( A1 => pipeline_stageD_target_Jump_temp_25_port, 
                           A2 => n17675, B1 => n17106, B2 => n15707, ZN => 
                           n15705);
   U10068 : AOI22_X1 port map( A1 => pipeline_data_to_RF_from_WB_25_port, A2 =>
                           n17332, B1 => pipeline_Alu_Out_Addr_to_mem_25_port, 
                           B2 => n17330, ZN => n15706);
   U9639 : AOI22_X1 port map( A1 => n17150, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N34, B1 => n17149,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_N66, ZN => 
                           n15196);
   U9638 : AOI22_X1 port map( A1 => n17359, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N164, B1 => n17126
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N132, ZN 
                           => n15197);
   U9637 : AOI22_X1 port map( A1 => n17419, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N229, B1 => n17681
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N261, ZN 
                           => n15198);
   U9636 : NAND4_X1 port map( A1 => n15196, A2 => n15197, A3 => n15198, A4 => 
                           n15199, ZN => n15195);
   U9635 : AOI211_X1 port map( C1 => n14993, C2 => n15014, A => n15194, B => 
                           n15195, ZN => n15193);
   U9634 : NAND2_X1 port map( A1 => n15192, A2 => n15193, ZN => 
                           pipeline_EXMEM_stage_N34);
   U9648 : AOI22_X1 port map( A1 => n17150, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N33, B1 => n17149,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_N65, ZN => 
                           n15210);
   U9647 : AOI22_X1 port map( A1 => n17359, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N163, B1 => n17126
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N131, ZN 
                           => n15211);
   U9646 : AOI22_X1 port map( A1 => n17419, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N228, B1 => n17681
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N260, ZN 
                           => n15212);
   U9645 : NAND4_X1 port map( A1 => n15210, A2 => n15211, A3 => n15212, A4 => 
                           n15213, ZN => n15209);
   U9644 : AOI211_X1 port map( C1 => n14993, C2 => n15015, A => n15208, B => 
                           n15209, ZN => n15207);
   U9643 : NAND2_X1 port map( A1 => n15206, A2 => n15207, ZN => 
                           pipeline_EXMEM_stage_N33);
   U10077 : AOI22_X1 port map( A1 => pipeline_stageF_PC_plus4_N31, A2 => n17108
                           , B1 => n17674, B2 => n13861, ZN => n15709);
   U10075 : AOI22_X1 port map( A1 => pipeline_stageD_target_Jump_temp_24_port, 
                           A2 => n17675, B1 => n17106, B2 => n15712, ZN => 
                           n15710);
   U10074 : AOI22_X1 port map( A1 => pipeline_data_to_RF_from_WB_24_port, A2 =>
                           n15605, B1 => pipeline_Alu_Out_Addr_to_mem_24_port, 
                           B2 => n17330, ZN => n15711);
   U9676 : AOI22_X1 port map( A1 => n17150, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N30, B1 => n17149,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_N62, ZN => 
                           n15255);
   U9880 : NOR2_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_2_port, A2 
                           => n15581, ZN => n14963);
   U9675 : AOI22_X1 port map( A1 => n14963, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N160, B1 => n17126
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N128, ZN 
                           => n15256);
   U9874 : NOR2_X1 port map( A1 => n17405, A2 => n15581, ZN => n14962);
   U9674 : AOI22_X1 port map( A1 => n14961, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N225, B1 => n14962
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N257, ZN 
                           => n15257);
   U9673 : NAND4_X1 port map( A1 => n15255, A2 => n15256, A3 => n15257, A4 => 
                           n15258, ZN => n15254);
   U9672 : AOI211_X1 port map( C1 => n14993, C2 => n15022, A => n15253, B => 
                           n15254, ZN => n15252);
   U9671 : NAND2_X1 port map( A1 => n15251, A2 => n15252, ZN => 
                           pipeline_EXMEM_stage_N30);
   U9660 : NOR2_X1 port map( A1 => n17159, A2 => n15224, ZN => n15225);
   U9658 : AOI22_X1 port map( A1 => n17150, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N32, B1 => n17149,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_N64, ZN => 
                           n15228);
   U9657 : AOI22_X1 port map( A1 => n17359, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N162, B1 => n14964
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N130, ZN 
                           => n15229);
   U9656 : AOI22_X1 port map( A1 => n14961, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N227, B1 => n17681
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N259, ZN 
                           => n15230);
   U9655 : AOI211_X1 port map( C1 => n14954, C2 => n15225, A => n15226, B => 
                           n15227, ZN => n15222);
   U9654 : OAI211_X1 port map( C1 => n15020, C2 => n14949, A => n15222, B => 
                           n15223, ZN => pipeline_EXMEM_stage_N32);
   U9723 : AOI22_X1 port map( A1 => n17150, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N26, B1 => n17149,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_N58, ZN => 
                           n15325);
   U9722 : AOI22_X1 port map( A1 => n14963, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N156, B1 => n17126
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N124, ZN 
                           => n15326);
   U9721 : AOI22_X1 port map( A1 => n14961, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N221, B1 => n14962
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N253, ZN 
                           => n15327);
   U9720 : NAND4_X1 port map( A1 => n15325, A2 => n15326, A3 => n15327, A4 => 
                           n15328, ZN => n15324);
   U9719 : AOI211_X1 port map( C1 => n14993, C2 => n15023, A => n15323, B => 
                           n15324, ZN => n15322);
   U9718 : NAND2_X1 port map( A1 => n15321, A2 => n15322, ZN => 
                           pipeline_EXMEM_stage_N26);
   U10083 : AOI22_X1 port map( A1 => pipeline_stageF_PC_plus4_N30, A2 => n17108
                           , B1 => n17674, B2 => n13860, ZN => n15714);
   U10081 : AOI22_X1 port map( A1 => pipeline_stageD_target_Jump_temp_23_port, 
                           A2 => n15607, B1 => n17106, B2 => n15717, ZN => 
                           n15715);
   U10080 : AOI22_X1 port map( A1 => pipeline_data_to_RF_from_WB_23_port, A2 =>
                           n15605, B1 => pipeline_Alu_Out_Addr_to_mem_23_port, 
                           B2 => n15606, ZN => n15716);
   U9709 : AOI22_X1 port map( A1 => n14965, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N27, B1 => n14966,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_N59, ZN => 
                           n15306);
   U9708 : AOI22_X1 port map( A1 => n14963, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N157, B1 => n17126
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N125, ZN 
                           => n15307);
   U9707 : AOI22_X1 port map( A1 => n17419, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N222, B1 => n14962
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N254, ZN 
                           => n15308);
   U9706 : NAND4_X1 port map( A1 => n15306, A2 => n15307, A3 => n15308, A4 => 
                           n15309, ZN => n15305);
   U9705 : AOI211_X1 port map( C1 => n14993, C2 => n15026, A => n15304, B => 
                           n15305, ZN => n15303);
   U9704 : NAND2_X1 port map( A1 => n15302, A2 => n15303, ZN => 
                           pipeline_EXMEM_stage_N27);
   U9700 : NOR2_X1 port map( A1 => pipeline_stageE_input1_to_ALU_21_port, A2 =>
                           n15285, ZN => n15286);
   U9697 : AOI22_X1 port map( A1 => n17150, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N28, B1 => n17149,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_N60, ZN => 
                           n15289);
   U9696 : AOI22_X1 port map( A1 => n14963, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N158, B1 => n17126
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N126, ZN 
                           => n15290);
   U9695 : AOI22_X1 port map( A1 => n14961, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N223, B1 => n14962
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N255, ZN 
                           => n15291);
   U9694 : AOI211_X1 port map( C1 => n17677, C2 => n15286, A => n15287, B => 
                           n15288, ZN => n15283);
   U9693 : OAI211_X1 port map( C1 => n15017, C2 => n14949, A => n15283, B => 
                           n15284, ZN => pipeline_EXMEM_stage_N28);
   U9793 : NOR2_X1 port map( A1 => pipeline_stageE_input1_to_ALU_11_port, A2 =>
                           n15449, ZN => n15450);
   U9791 : AOI22_X1 port map( A1 => n17150, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N18, B1 => n17149,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_N50, ZN => 
                           n15453);
   U9790 : AOI22_X1 port map( A1 => n17680, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N148, B1 => n17126
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N116, ZN 
                           => n15454);
   U9789 : AOI22_X1 port map( A1 => n17419, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N213, B1 => n17360
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N245, ZN 
                           => n15455);
   U9788 : AOI211_X1 port map( C1 => n17677, C2 => n15450, A => n15451, B => 
                           n15452, ZN => n15447);
   U9787 : OAI211_X1 port map( C1 => n15040, C2 => n14949, A => n15447, B => 
                           n15448, ZN => pipeline_EXMEM_stage_N18);
   U9784 : NOR2_X1 port map( A1 => pipeline_stageE_input1_to_ALU_12_port, A2 =>
                           n15435, ZN => n15436);
   U9783 : AOI22_X1 port map( A1 => n17150, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N19, B1 => n17149,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_N51, ZN => 
                           n15439);
   U9782 : AOI22_X1 port map( A1 => n17680, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N149, B1 => n17126
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N117, ZN 
                           => n15440);
   U9781 : AOI22_X1 port map( A1 => n14961, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N214, B1 => n17360
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N246, ZN 
                           => n15441);
   U9780 : AOI211_X1 port map( C1 => n17677, C2 => n15436, A => n15437, B => 
                           n15438, ZN => n15433);
   U9779 : OAI211_X1 port map( C1 => n15030, C2 => n14949, A => n15433, B => 
                           n15434, ZN => pipeline_EXMEM_stage_N19);
   U9731 : AOI22_X1 port map( A1 => n17150, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N25, B1 => n17149,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_N57, ZN => 
                           n15340);
   U9730 : AOI22_X1 port map( A1 => n17680, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N155, B1 => n17126
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N123, ZN 
                           => n15341);
   U9729 : AOI22_X1 port map( A1 => n14961, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N220, B1 => n17360
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N252, ZN 
                           => n15342);
   U9728 : NAND4_X1 port map( A1 => n15340, A2 => n15341, A3 => n15342, A4 => 
                           n15343, ZN => n15339);
   U9727 : AOI211_X1 port map( C1 => n14993, C2 => n15021, A => n15338, B => 
                           n15339, ZN => n15337);
   U9726 : NAND2_X1 port map( A1 => n15336, A2 => n15337, ZN => 
                           pipeline_EXMEM_stage_N25);
   U9775 : AOI22_X1 port map( A1 => n17150, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N20, B1 => n17149,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_N52, ZN => 
                           n15421);
   U9774 : AOI22_X1 port map( A1 => n17680, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N150, B1 => n17126
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N118, ZN 
                           => n15422);
   U9773 : AOI22_X1 port map( A1 => n14961, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N215, B1 => n14962
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N247, ZN 
                           => n15423);
   U9772 : NAND4_X1 port map( A1 => n15421, A2 => n15422, A3 => n15423, A4 => 
                           n15424, ZN => n15420);
   U9771 : AOI211_X1 port map( C1 => n14993, C2 => n15033, A => n15419, B => 
                           n15420, ZN => n15418);
   U9770 : NAND2_X1 port map( A1 => n15417, A2 => n15418, ZN => 
                           pipeline_EXMEM_stage_N20);
   U9760 : NOR2_X1 port map( A1 => pipeline_stageE_input1_to_ALU_15_port, A2 =>
                           n15386, ZN => n15387);
   U9758 : AOI22_X1 port map( A1 => n17150, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N22, B1 => n17149,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_N54, ZN => 
                           n15390);
   U9757 : AOI22_X1 port map( A1 => n14963, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N152, B1 => n17126
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N120, ZN 
                           => n15391);
   U9756 : AOI22_X1 port map( A1 => n14961, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N217, B1 => n14962
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N249, ZN 
                           => n15392);
   U9755 : AOI211_X1 port map( C1 => n17677, C2 => n15387, A => n15388, B => 
                           n15389, ZN => n15384);
   U9754 : OAI211_X1 port map( C1 => n15029, C2 => n14949, A => n15384, B => 
                           n15385, ZN => pipeline_EXMEM_stage_N22);
   U9669 : AOI22_X1 port map( A1 => n14965, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N31, B1 => n17149,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_N63, ZN => 
                           n15240);
   U9668 : AOI22_X1 port map( A1 => n14963, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N161, B1 => n17126
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N129, ZN 
                           => n15241);
   U9667 : AOI22_X1 port map( A1 => n14961, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N226, B1 => n17681
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N258, ZN 
                           => n15242);
   U9666 : NAND4_X1 port map( A1 => n15240, A2 => n15241, A3 => n15242, A4 => 
                           n15243, ZN => n15239);
   U9665 : AOI211_X1 port map( C1 => n14993, C2 => n15013, A => n15238, B => 
                           n15239, ZN => n15237);
   U9664 : NAND2_X1 port map( A1 => n15236, A2 => n15237, ZN => 
                           pipeline_EXMEM_stage_N31);
   U9868 : NAND2_X1 port map( A1 => pipeline_stageE_input1_to_ALU_4_port, A2 =>
                           n14952, ZN => n15556);
   U9865 : AOI22_X1 port map( A1 => n17150, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N11, B1 => n17149,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_N43, ZN => 
                           n15560);
   U9864 : AOI22_X1 port map( A1 => n17359, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N141, B1 => n17126
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N109, ZN 
                           => n15561);
   U9863 : AOI22_X1 port map( A1 => n17419, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N206, B1 => n17681
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N238, ZN 
                           => n15562);
   U9862 : NAND4_X1 port map( A1 => n15560, A2 => n15561, A3 => n15562, A4 => 
                           n15563, ZN => n15559);
   U9861 : AOI211_X1 port map( C1 => n14993, C2 => n15041, A => n15558, B => 
                           n15559, ZN => n15557);
   U9860 : OAI21_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, B2 
                           => n15556, A => n15557, ZN => 
                           pipeline_EXMEM_stage_N11);
   U10089 : AOI22_X1 port map( A1 => pipeline_stageF_PC_plus4_N29, A2 => n15610
                           , B1 => n17674, B2 => n13859, ZN => n15719);
   U10087 : AOI22_X1 port map( A1 => pipeline_stageD_target_Jump_temp_22_port, 
                           A2 => n17676, B1 => n17106, B2 => n15722, ZN => 
                           n15720);
   U10086 : AOI22_X1 port map( A1 => pipeline_data_to_RF_from_WB_22_port, A2 =>
                           n15605, B1 => pipeline_Alu_Out_Addr_to_mem_22_port, 
                           B2 => n15606, ZN => n15721);
   U9854 : AOI22_X1 port map( A1 => n17150, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N12, B1 => n17149,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_N44, ZN => 
                           n15547);
   U9853 : AOI22_X1 port map( A1 => n17359, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N142, B1 => n17126
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N110, ZN 
                           => n15548);
   U9852 : AOI22_X1 port map( A1 => n17419, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N207, B1 => n17681
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N239, ZN 
                           => n15549);
   U9851 : NAND4_X1 port map( A1 => n15547, A2 => n15548, A3 => n15549, A4 => 
                           n15550, ZN => n15546);
   U9850 : AOI211_X1 port map( C1 => n14993, C2 => n15042, A => n15545, B => 
                           n15546, ZN => n15544);
   U9849 : NAND2_X1 port map( A1 => n15543, A2 => n15544, ZN => 
                           pipeline_EXMEM_stage_N12);
   U9844 : AOI22_X1 port map( A1 => n14965, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N13, B1 => n17149,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_N45, ZN => 
                           n15532);
   U9843 : AOI22_X1 port map( A1 => n17359, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N143, B1 => n17126
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N111, ZN 
                           => n15533);
   U9842 : AOI22_X1 port map( A1 => n17419, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N208, B1 => n17681
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N240, ZN 
                           => n15534);
   U9841 : NAND4_X1 port map( A1 => n15532, A2 => n15533, A3 => n15534, A4 => 
                           n15535, ZN => n15531);
   U9840 : AOI211_X1 port map( C1 => n14993, C2 => n15043, A => n15530, B => 
                           n15531, ZN => n15529);
   U9839 : NAND2_X1 port map( A1 => n15528, A2 => n15529, ZN => 
                           pipeline_EXMEM_stage_N13);
   U9465 : NOR2_X1 port map( A1 => n12649, A2 => n17740, ZN => n14955);
   U9463 : AOI22_X1 port map( A1 => n17150, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N9, B1 => n17149, 
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_N41, ZN => 
                           n14958);
   U9462 : AOI22_X1 port map( A1 => n17680, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N139, B1 => n17126
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N107, ZN 
                           => n14959);
   U9461 : AOI22_X1 port map( A1 => n17419, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N204, B1 => n17360
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N236, ZN 
                           => n14960);
   U9460 : AOI211_X1 port map( C1 => n14954, C2 => n14955, A => n14956, B => 
                           n14957, ZN => n14950);
   U9459 : OAI211_X1 port map( C1 => n14948, C2 => n14949, A => n14950, B => 
                           n14951, ZN => pipeline_EXMEM_stage_N9);
   U9890 : NOR2_X1 port map( A1 => n17739, A2 => 
                           pipeline_stageE_input1_to_ALU_3_port, ZN => n15574);
   U9883 : AOI22_X1 port map( A1 => n17150, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N10, B1 => n14966,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_N42, ZN => 
                           n15577);
   U9877 : AOI22_X1 port map( A1 => n17359, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N140, B1 => n14964
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N108, ZN 
                           => n15578);
   U9873 : AOI22_X1 port map( A1 => n17419, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N205, B1 => n17681
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N237, ZN 
                           => n15579);
   U9872 : AOI211_X1 port map( C1 => n17677, C2 => n15574, A => n15575, B => 
                           n15576, ZN => n15570);
   U9869 : OAI211_X1 port map( C1 => n15045, C2 => n14949, A => n15570, B => 
                           n15571, ZN => pipeline_EXMEM_stage_N10);
   U9688 : AOI22_X1 port map( A1 => n17150, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N29, B1 => n17149,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_N61, ZN => 
                           n15273);
   U9687 : AOI22_X1 port map( A1 => n14963, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N159, B1 => n17126
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N127, ZN 
                           => n15274);
   U9686 : AOI22_X1 port map( A1 => n14961, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N224, B1 => n14962
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N256, ZN 
                           => n15275);
   U9685 : NAND4_X1 port map( A1 => n15273, A2 => n15274, A3 => n15275, A4 => 
                           n15276, ZN => n15272);
   U9684 : AOI211_X1 port map( C1 => n14993, C2 => n15024, A => n15271, B => 
                           n15272, ZN => n15270);
   U9683 : NAND2_X1 port map( A1 => n15269, A2 => n15270, ZN => 
                           pipeline_EXMEM_stage_N29);
   U9470 : AOI22_X1 port map( A1 => n17150, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N8, B1 => n17149, 
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_N40, ZN => 
                           n14977);
   U9469 : AOI22_X1 port map( A1 => n17680, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N138, B1 => n17126
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N106, ZN 
                           => n14978);
   U9468 : AOI22_X1 port map( A1 => n17419, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N203, B1 => n17360
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N235, ZN 
                           => n14979);
   U9467 : NOR3_X1 port map( A1 => n14974, A2 => n14975, A3 => n14976, ZN => 
                           n14971);
   U9466 : OAI211_X1 port map( C1 => n14970, C2 => n14949, A => n14971, B => 
                           n14972, ZN => pipeline_EXMEM_stage_N8);
   U9742 : AOI22_X1 port map( A1 => n17150, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N24, B1 => n17149,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_N56, ZN => 
                           n15357);
   U9741 : AOI22_X1 port map( A1 => n17680, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N154, B1 => n17126
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N122, ZN 
                           => n15358);
   U9740 : AOI22_X1 port map( A1 => n14961, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N219, B1 => n17360
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N251, ZN 
                           => n15359);
   U9739 : NAND4_X1 port map( A1 => n15357, A2 => n15358, A3 => n15359, A4 => 
                           n15360, ZN => n15356);
   U9738 : AOI211_X1 port map( C1 => n14993, C2 => n15025, A => n15355, B => 
                           n15356, ZN => n15354);
   U9737 : NAND2_X1 port map( A1 => n15353, A2 => n15354, ZN => 
                           pipeline_EXMEM_stage_N24);
   U9752 : NOR2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_A_16_port, A2 
                           => n15372, ZN => n15373);
   U9750 : AOI22_X1 port map( A1 => n17150, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N23, B1 => n14966,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_N55, ZN => 
                           n15376);
   U9749 : AOI22_X1 port map( A1 => n14963, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N153, B1 => n14964
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N121, ZN 
                           => n15377);
   U9748 : AOI22_X1 port map( A1 => n14961, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N218, B1 => n17681
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N250, ZN 
                           => n15378);
   U9747 : AOI211_X1 port map( C1 => n17677, C2 => n15373, A => n15374, B => 
                           n15375, ZN => n15370);
   U9746 : OAI211_X1 port map( C1 => n15032, C2 => n14949, A => n15370, B => 
                           n15371, ZN => pipeline_EXMEM_stage_N23);
   U9825 : NOR2_X1 port map( A1 => pipeline_stageE_input1_to_ALU_8_port, A2 => 
                           n15498, ZN => n15499);
   U9823 : AOI22_X1 port map( A1 => n17150, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N15, B1 => n17149,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_N47, ZN => 
                           n15502);
   U9822 : AOI22_X1 port map( A1 => n17359, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N145, B1 => n17126
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N113, ZN 
                           => n15503);
   U9821 : AOI22_X1 port map( A1 => n17419, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N210, B1 => n17360
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N242, ZN 
                           => n15504);
   U9820 : AOI211_X1 port map( C1 => n17677, C2 => n15499, A => n15500, B => 
                           n15501, ZN => n15496);
   U9819 : OAI211_X1 port map( C1 => n15039, C2 => n14949, A => n15496, B => 
                           n15497, ZN => pipeline_EXMEM_stage_N15);
   U9803 : AOI22_X1 port map( A1 => n17150, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N17, B1 => n17149,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_N49, ZN => 
                           n15468);
   U9802 : AOI22_X1 port map( A1 => n17680, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N147, B1 => n17126
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N115, ZN 
                           => n15469);
   U9801 : AOI22_X1 port map( A1 => n17419, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N212, B1 => n17360
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N244, ZN 
                           => n15470);
   U9800 : NAND4_X1 port map( A1 => n15468, A2 => n15469, A3 => n15470, A4 => 
                           n15471, ZN => n15467);
   U9799 : AOI211_X1 port map( C1 => n14993, C2 => n15034, A => n15466, B => 
                           n15467, ZN => n15465);
   U9798 : NAND2_X1 port map( A1 => n15464, A2 => n15465, ZN => 
                           pipeline_EXMEM_stage_N17);
   U9815 : AOI22_X1 port map( A1 => n17150, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N16, B1 => n17149,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_N48, ZN => 
                           n15486);
   U9814 : AOI22_X1 port map( A1 => n17680, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N146, B1 => n17126
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N114, ZN 
                           => n15487);
   U9813 : AOI22_X1 port map( A1 => n17419, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N211, B1 => n17360
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N243, ZN 
                           => n15488);
   U9812 : NAND4_X1 port map( A1 => n15486, A2 => n15487, A3 => n15488, A4 => 
                           n15489, ZN => n15485);
   U9811 : AOI211_X1 port map( C1 => n14993, C2 => n15035, A => n15484, B => 
                           n15485, ZN => n15483);
   U9810 : NAND2_X1 port map( A1 => n15482, A2 => n15483, ZN => 
                           pipeline_EXMEM_stage_N16);
   U9833 : NOR2_X1 port map( A1 => pipeline_stageE_input1_to_ALU_7_port, A2 => 
                           n15512, ZN => n15513);
   U9831 : AOI22_X1 port map( A1 => n17150, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N14, B1 => n17149,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_N46, ZN => 
                           n15516);
   U9830 : AOI22_X1 port map( A1 => n17359, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N144, B1 => n14964
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N112, ZN 
                           => n15517);
   U9829 : AOI22_X1 port map( A1 => n17419, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N209, B1 => n17360
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N241, ZN 
                           => n15518);
   U9828 : AOI211_X1 port map( C1 => n17677, C2 => n15513, A => n15514, B => 
                           n15515, ZN => n15510);
   U9827 : OAI211_X1 port map( C1 => n15037, C2 => n14949, A => n15510, B => 
                           n15511, ZN => pipeline_EXMEM_stage_N14);
   U9767 : AOI22_X1 port map( A1 => n17150, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N21, B1 => n17149,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_N53, ZN => 
                           n15405);
   U9766 : AOI22_X1 port map( A1 => n17680, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N151, B1 => n17126
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N119, ZN 
                           => n15406);
   U9765 : AOI22_X1 port map( A1 => n14961, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N216, B1 => n14962
                           , B2 => pipeline_stageE_EXE_ALU_alu_shift_N248, ZN 
                           => n15407);
   U9764 : NAND4_X1 port map( A1 => n15405, A2 => n15406, A3 => n15407, A4 => 
                           n15408, ZN => n15404);
   U9763 : AOI211_X1 port map( C1 => n14993, C2 => n15027, A => n15403, B => 
                           n15404, ZN => n15402);
   U9762 : NAND2_X1 port map( A1 => n15401, A2 => n15402, ZN => 
                           pipeline_EXMEM_stage_N21);
   U10095 : AOI22_X1 port map( A1 => pipeline_stageF_PC_plus4_N28, A2 => n15610
                           , B1 => n17674, B2 => n13858, ZN => n15724);
   U10093 : AOI22_X1 port map( A1 => pipeline_stageD_target_Jump_temp_21_port, 
                           A2 => n17675, B1 => n15608, B2 => n15727, ZN => 
                           n15725);
   U10092 : AOI22_X1 port map( A1 => pipeline_data_to_RF_from_WB_21_port, A2 =>
                           n15605, B1 => pipeline_Alu_Out_Addr_to_mem_21_port, 
                           B2 => n15606, ZN => n15726);
   U9981 : AOI22_X1 port map( A1 => pipeline_inst_IFID_DEC_31_port, A2 => 
                           n15600, B1 => n17673, B2 => InstrFetched_31_port, ZN
                           => n15653);
   U9973 : AOI22_X1 port map( A1 => pipeline_inst_IFID_DEC_27_port, A2 => 
                           n15600, B1 => n17107, B2 => InstrFetched_27_port, ZN
                           => n15649);
   U9969 : AOI22_X1 port map( A1 => 
                           pipeline_stageD_offset_jump_sign_ext_31_port, A2 => 
                           n15600, B1 => n17107, B2 => InstrFetched_25_port, ZN
                           => n15645);
   U9961 : AOI22_X1 port map( A1 => 
                           pipeline_stageD_offset_jump_sign_ext_21_port, A2 => 
                           n17671, B1 => n17107, B2 => InstrFetched_21_port, ZN
                           => n15641);
   U9977 : AOI22_X1 port map( A1 => pipeline_inst_IFID_DEC_29_port, A2 => 
                           n15600, B1 => n17673, B2 => InstrFetched_29_port, ZN
                           => n15651);
   U9963 : AOI22_X1 port map( A1 => 
                           pipeline_stageD_offset_jump_sign_ext_22_port, A2 => 
                           n15600, B1 => n17107, B2 => InstrFetched_22_port, ZN
                           => n15642);
   U10145 : AOI22_X1 port map( A1 => n15600, A2 => 
                           pipeline_nextPC_IFID_DEC_8_port, B1 => n17673, B2 =>
                           pipeline_stageF_PC_plus4_N15, ZN => n15768);
   U10156 : AOI22_X1 port map( A1 => n15600, A2 => 
                           pipeline_nextPC_IFID_DEC_3_port, B1 => n17673, B2 =>
                           pipeline_stageF_PC_plus4_N10, ZN => n15778);
   U10067 : AOI22_X1 port map( A1 => n15600, A2 => 
                           pipeline_nextPC_IFID_DEC_26_port, B1 => n17673, B2 
                           => pipeline_stageF_PC_plus4_N33, ZN => n15703);
   U9941 : AOI22_X1 port map( A1 => n15600, A2 => 
                           pipeline_stageD_offset_to_jump_temp_10_port, B1 => 
                           n17673, B2 => InstrFetched_10_port, ZN => n15631);
   U9965 : AOI22_X1 port map( A1 => 
                           pipeline_stageD_offset_jump_sign_ext_23_port, A2 => 
                           n17671, B1 => n17107, B2 => InstrFetched_23_port, ZN
                           => n15643);
   U10055 : AOI22_X1 port map( A1 => n15600, A2 => 
                           pipeline_nextPC_IFID_DEC_28_port, B1 => n15601, B2 
                           => pipeline_stageF_PC_plus4_N35, ZN => n15693);
   U10198 : AOI22_X1 port map( A1 => n17671, A2 => 
                           pipeline_nextPC_IFID_DEC_10_port, B1 => n17107, B2 
                           => pipeline_stageF_PC_plus4_N17, ZN => n15813);
   U10174 : AOI22_X1 port map( A1 => n15600, A2 => 
                           pipeline_nextPC_IFID_DEC_5_port, B1 => n15601, B2 =>
                           pipeline_stageF_PC_plus4_N12, ZN => n15793);
   U9931 : AOI22_X1 port map( A1 => n17671, A2 => 
                           pipeline_stageD_offset_to_jump_temp_5_port, B1 => 
                           n17107, B2 => InstrFetched_5_port, ZN => n15626);
   U10091 : AOI22_X1 port map( A1 => n15600, A2 => 
                           pipeline_nextPC_IFID_DEC_22_port, B1 => n17107, B2 
                           => pipeline_stageF_PC_plus4_N29, ZN => n15723);
   U10109 : AOI22_X1 port map( A1 => n15600, A2 => 
                           pipeline_nextPC_IFID_DEC_19_port, B1 => n17107, B2 
                           => pipeline_stageF_PC_plus4_N26, ZN => n15738);
   U9953 : AOI22_X1 port map( A1 => n15600, A2 => 
                           pipeline_stageD_offset_jump_sign_ext_17_port, B1 => 
                           n15601, B2 => InstrFetched_17_port, ZN => n15637);
   U10168 : AOI22_X1 port map( A1 => n15600, A2 => 
                           pipeline_nextPC_IFID_DEC_4_port, B1 => n15601, B2 =>
                           pipeline_stageF_PC_plus4_N11, ZN => n15788);
   U9929 : AOI22_X1 port map( A1 => n17671, A2 => 
                           pipeline_stageD_offset_to_jump_temp_4_port, B1 => 
                           n17107, B2 => InstrFetched_4_port, ZN => n15625);
   U10079 : AOI22_X1 port map( A1 => n17671, A2 => 
                           pipeline_nextPC_IFID_DEC_24_port, B1 => n17673, B2 
                           => pipeline_stageF_PC_plus4_N31, ZN => n15713);
   U10139 : AOI22_X1 port map( A1 => n17671, A2 => 
                           pipeline_nextPC_IFID_DEC_13_port, B1 => n17673, B2 
                           => pipeline_stageF_PC_plus4_N20, ZN => n15763);
   U9905 : AOI22_X1 port map( A1 => n17671, A2 => 
                           pipeline_stageD_offset_to_jump_temp_14_port, B1 => 
                           n17673, B2 => InstrFetched_14_port, ZN => n15599);
   U9951 : AOI22_X1 port map( A1 => n17671, A2 => 
                           pipeline_stageD_offset_jump_sign_ext_16_port, B1 => 
                           n17673, B2 => InstrFetched_16_port, ZN => n15636);
   U10162 : AOI22_X1 port map( A1 => n17671, A2 => 
                           pipeline_nextPC_IFID_DEC_7_port, B1 => n17673, B2 =>
                           pipeline_stageF_PC_plus4_N14, ZN => n15783);
   U10230 : AOI22_X1 port map( A1 => n17671, A2 => 
                           pipeline_nextPC_IFID_DEC_30_port, B1 => n17107, B2 
                           => pipeline_stageF_PC_plus4_N37, ZN => n15837);
   U9957 : AOI22_X1 port map( A1 => n17671, A2 => 
                           pipeline_stageD_offset_jump_sign_ext_19_port, B1 => 
                           n17107, B2 => InstrFetched_19_port, ZN => n15639);
   U10210 : AOI22_X1 port map( A1 => n17671, A2 => 
                           pipeline_nextPC_IFID_DEC_2_port, B1 => n17107, B2 =>
                           pipeline_stageF_PC_plus4_N9, ZN => n15823);
   U9959 : AOI22_X1 port map( A1 => n17671, A2 => 
                           pipeline_stageD_offset_jump_sign_ext_20_port, B1 => 
                           n17107, B2 => InstrFetched_20_port, ZN => n15640);
   U10127 : AOI22_X1 port map( A1 => n17671, A2 => 
                           pipeline_nextPC_IFID_DEC_15_port, B1 => n17107, B2 
                           => pipeline_stageF_PC_plus4_N22, ZN => n15753);
   U10121 : AOI22_X1 port map( A1 => n17671, A2 => 
                           pipeline_nextPC_IFID_DEC_17_port, B1 => n17672, B2 
                           => pipeline_stageF_PC_plus4_N24, ZN => n15748);
   U10103 : AOI22_X1 port map( A1 => n17671, A2 => 
                           pipeline_nextPC_IFID_DEC_20_port, B1 => n17107, B2 
                           => pipeline_stageF_PC_plus4_N27, ZN => n15733);
   U9939 : AOI22_X1 port map( A1 => n17671, A2 => 
                           pipeline_stageD_offset_to_jump_temp_9_port, B1 => 
                           n17107, B2 => InstrFetched_9_port, ZN => n15630);
   U9947 : AOI22_X1 port map( A1 => n15600, A2 => 
                           pipeline_stageD_offset_to_jump_temp_13_port, B1 => 
                           n17673, B2 => InstrFetched_13_port, ZN => n15634);
   U9943 : AOI22_X1 port map( A1 => n15600, A2 => 
                           pipeline_stageD_offset_to_jump_temp_11_port, B1 => 
                           n17673, B2 => InstrFetched_11_port, ZN => n15632);
   U10073 : AOI22_X1 port map( A1 => n15600, A2 => 
                           pipeline_nextPC_IFID_DEC_25_port, B1 => n17673, B2 
                           => pipeline_stageF_PC_plus4_N32, ZN => n15708);
   U10097 : AOI22_X1 port map( A1 => n15600, A2 => 
                           pipeline_nextPC_IFID_DEC_21_port, B1 => n17672, B2 
                           => pipeline_stageF_PC_plus4_N28, ZN => n15728);
   U9923 : AOI22_X1 port map( A1 => n17671, A2 => 
                           pipeline_stageD_offset_to_jump_temp_1_port, B1 => 
                           n15601, B2 => InstrFetched_1_port, ZN => n15622);
   U9933 : AOI22_X1 port map( A1 => n17671, A2 => 
                           pipeline_stageD_offset_to_jump_temp_6_port, B1 => 
                           n17107, B2 => InstrFetched_6_port, ZN => n15627);
   U9945 : AOI22_X1 port map( A1 => n15600, A2 => 
                           pipeline_stageD_offset_to_jump_temp_12_port, B1 => 
                           n15601, B2 => InstrFetched_12_port, ZN => n15633);
   U10061 : AOI22_X1 port map( A1 => n15600, A2 => 
                           pipeline_nextPC_IFID_DEC_27_port, B1 => n15601, B2 
                           => pipeline_stageF_PC_plus4_N34, ZN => n15698);
   U10204 : AOI22_X1 port map( A1 => n17671, A2 => 
                           pipeline_nextPC_IFID_DEC_12_port, B1 => n17107, B2 
                           => pipeline_stageF_PC_plus4_N19, ZN => n15818);
   U10192 : AOI22_X1 port map( A1 => n17671, A2 => 
                           pipeline_nextPC_IFID_DEC_9_port, B1 => n17672, B2 =>
                           pipeline_stageF_PC_plus4_N16, ZN => n15808);
   U10186 : AOI22_X1 port map( A1 => n15600, A2 => 
                           pipeline_nextPC_IFID_DEC_11_port, B1 => n17107, B2 
                           => pipeline_stageF_PC_plus4_N18, ZN => n15803);
   U10226 : AOI22_X1 port map( A1 => n15600, A2 => 
                           pipeline_nextPC_IFID_DEC_1_port, B1 => n17107, B2 =>
                           pipeline_stageF_PC_plus4_N8, ZN => n15835);
   U9955 : AOI22_X1 port map( A1 => n15600, A2 => 
                           pipeline_stageD_offset_jump_sign_ext_18_port, B1 => 
                           n17673, B2 => InstrFetched_18_port, ZN => n15638);
   U9949 : AOI22_X1 port map( A1 => n15600, A2 => 
                           pipeline_stageD_offset_to_jump_temp_15_port, B1 => 
                           n17673, B2 => InstrFetched_15_port, ZN => n15635);
   U10101 : AOI22_X1 port map( A1 => pipeline_stageF_PC_plus4_N27, A2 => n15610
                           , B1 => n17674, B2 => n13857, ZN => n15729);
   U10099 : AOI22_X1 port map( A1 => pipeline_stageD_target_Jump_temp_20_port, 
                           A2 => n15607, B1 => n17106, B2 => n15732, ZN => 
                           n15730);
   U10098 : AOI22_X1 port map( A1 => pipeline_data_to_RF_from_WB_20_port, A2 =>
                           n15605, B1 => pipeline_Alu_Out_Addr_to_mem_20_port, 
                           B2 => n15606, ZN => n15731);
   U10202 : AOI22_X1 port map( A1 => pipeline_stageF_PC_plus4_N19, A2 => n17108
                           , B1 => n17674, B2 => n13813, ZN => n15814);
   U10200 : AOI22_X1 port map( A1 => pipeline_stageD_target_Jump_temp_12_port, 
                           A2 => n17675, B1 => n17106, B2 => n15817, ZN => 
                           n15815);
   U10199 : AOI22_X1 port map( A1 => pipeline_data_to_RF_from_WB_12_port, A2 =>
                           n17332, B1 => pipeline_Alu_Out_Addr_to_mem_12_port, 
                           B2 => n17330, ZN => n15816);
   U10143 : AOI22_X1 port map( A1 => pipeline_stageF_PC_plus4_N15, A2 => n17108
                           , B1 => n17674, B2 => n13850, ZN => n15764);
   U10141 : AOI22_X1 port map( A1 => pipeline_stageD_target_Jump_temp_8_port, 
                           A2 => n17676, B1 => n17106, B2 => n15767, ZN => 
                           n15765);
   U10140 : AOI22_X1 port map( A1 => pipeline_data_to_RF_from_WB_8_port, A2 => 
                           n17333, B1 => pipeline_Alu_Out_Addr_to_mem_8_port, 
                           B2 => n15606, ZN => n15766);
   U10113 : AOI22_X1 port map( A1 => pipeline_stageF_PC_plus4_N25, A2 => n17108
                           , B1 => n17674, B2 => n13855, ZN => n15739);
   U10111 : AOI22_X1 port map( A1 => pipeline_stageD_target_Jump_temp_18_port, 
                           A2 => n17675, B1 => n17106, B2 => n15742, ZN => 
                           n15740);
   U10110 : AOI22_X1 port map( A1 => pipeline_data_to_RF_from_WB_18_port, A2 =>
                           n15605, B1 => pipeline_Alu_Out_Addr_to_mem_18_port, 
                           B2 => n15606, ZN => n15741);
   U10125 : AOI22_X1 port map( A1 => pipeline_stageF_PC_plus4_N22, A2 => n17108
                           , B1 => n15611, B2 => n13853, ZN => n15749);
   U10123 : AOI22_X1 port map( A1 => pipeline_stageD_target_Jump_temp_15_port, 
                           A2 => n17676, B1 => n17106, B2 => n15752, ZN => 
                           n15750);
   U10122 : AOI22_X1 port map( A1 => pipeline_data_to_RF_from_WB_15_port, A2 =>
                           n17333, B1 => pipeline_Alu_Out_Addr_to_mem_15_port, 
                           B2 => n17331, ZN => n15751);
   U10154 : AOI22_X1 port map( A1 => pipeline_stageF_PC_plus4_N10, A2 => n17108
                           , B1 => n15611, B2 => n13845, ZN => n15774);
   U10152 : AOI22_X1 port map( A1 => pipeline_stageD_target_Jump_temp_3_port, 
                           A2 => n15607, B1 => n17106, B2 => n15777, ZN => 
                           n15775);
   U10151 : AOI22_X1 port map( A1 => pipeline_Alu_Out_Addr_to_mem_3_port, A2 =>
                           n17330, B1 => pipeline_data_to_RF_from_WB_3_port, B2
                           => n17333, ZN => n15776);
   U9909 : AOI22_X1 port map( A1 => pipeline_stageF_PC_plus4_N23, A2 => n17108,
                           B1 => n17674, B2 => n13945, ZN => n15602);
   U9907 : AOI22_X1 port map( A1 => pipeline_stageD_target_Jump_temp_16_port, 
                           A2 => n17676, B1 => n17106, B2 => n15609, ZN => 
                           n15603);
   U9906 : AOI22_X1 port map( A1 => pipeline_data_to_RF_from_WB_16_port, A2 => 
                           n17333, B1 => pipeline_Alu_Out_Addr_to_mem_16_port, 
                           B2 => n17331, ZN => n15604);
   U10196 : AOI22_X1 port map( A1 => pipeline_stageF_PC_plus4_N17, A2 => n15610
                           , B1 => n17674, B2 => n13817, ZN => n15809);
   U10194 : AOI22_X1 port map( A1 => pipeline_stageD_target_Jump_temp_10_port, 
                           A2 => n17676, B1 => n17106, B2 => n15812, ZN => 
                           n15810);
   U10193 : AOI22_X1 port map( A1 => pipeline_data_to_RF_from_WB_10_port, A2 =>
                           n17332, B1 => pipeline_Alu_Out_Addr_to_mem_10_port, 
                           B2 => n17330, ZN => n15811);
   U10166 : AOI22_X1 port map( A1 => pipeline_stageF_PC_plus4_N11, A2 => n17108
                           , B1 => n15611, B2 => n13837, ZN => n15784);
   U10164 : AOI22_X1 port map( A1 => pipeline_stageD_target_Jump_temp_4_port, 
                           A2 => n17675, B1 => n17106, B2 => n15787, ZN => 
                           n15785);
   U10163 : AOI22_X1 port map( A1 => pipeline_data_to_RF_from_WB_4_port, A2 => 
                           n17333, B1 => pipeline_Alu_Out_Addr_to_mem_4_port, 
                           B2 => n17331, ZN => n15786);
   U10208 : AOI22_X1 port map( A1 => pipeline_stageF_PC_plus4_N9, A2 => n17108,
                           B1 => n15611, B2 => n13810, ZN => n15819);
   U10206 : AOI22_X1 port map( A1 => pipeline_stageD_target_Jump_temp_2_port, 
                           A2 => n15607, B1 => n17106, B2 => n15822, ZN => 
                           n15820);
   U10205 : AOI22_X1 port map( A1 => pipeline_data_to_RF_from_WB_2_port, A2 => 
                           n17332, B1 => pipeline_Alu_Out_Addr_to_mem_2_port, 
                           B2 => n17330, ZN => n15821);
   U10133 : AOI22_X1 port map( A1 => n15600, A2 => 
                           pipeline_nextPC_IFID_DEC_14_port, B1 => n17107, B2 
                           => pipeline_stageF_PC_plus4_N21, ZN => n15758);
   U10115 : AOI22_X1 port map( A1 => n15600, A2 => 
                           pipeline_nextPC_IFID_DEC_18_port, B1 => n17107, B2 
                           => pipeline_stageF_PC_plus4_N25, ZN => n15743);
   U9937 : AOI22_X1 port map( A1 => n15600, A2 => 
                           pipeline_stageD_offset_to_jump_temp_8_port, B1 => 
                           n17107, B2 => InstrFetched_8_port, ZN => n15629);
   U10228 : AOI22_X1 port map( A1 => n15600, A2 => 
                           pipeline_nextPC_IFID_DEC_29_port, B1 => n17107, B2 
                           => pipeline_stageF_PC_plus4_N36, ZN => n15836);
   U10048 : AOI222_X1 port map( A1 => n17331, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_31_port, B1 => 
                           pipeline_stageD_target_Jump_temp_31_port, B2 => 
                           n17675, C1 => n17106, C2 => n15688, ZN => n15686);
   U10047 : AOI22_X1 port map( A1 => pipeline_data_to_RF_from_WB_31_port, A2 =>
                           n17332, B1 => n17674, B2 => n13938, ZN => n15687);
   U10046 : NAND2_X1 port map( A1 => n15686, A2 => n15687, ZN => n3924);
   U10178 : AOI22_X1 port map( A1 => pipeline_stageF_PC_plus4_N13, A2 => n17108
                           , B1 => n15611, B2 => n13829, ZN => n15794);
   U10176 : AOI22_X1 port map( A1 => pipeline_stageD_target_Jump_temp_6_port, 
                           A2 => n17676, B1 => n17106, B2 => n15797, ZN => 
                           n15795);
   U10175 : AOI22_X1 port map( A1 => pipeline_data_to_RF_from_WB_6_port, A2 => 
                           n17333, B1 => pipeline_Alu_Out_Addr_to_mem_6_port, 
                           B2 => n17331, ZN => n15796);
   U10137 : AOI22_X1 port map( A1 => pipeline_stageF_PC_plus4_N20, A2 => n17108
                           , B1 => n17674, B2 => n13851, ZN => n15759);
   U10135 : AOI22_X1 port map( A1 => pipeline_stageD_target_Jump_temp_13_port, 
                           A2 => n15607, B1 => n17106, B2 => n15762, ZN => 
                           n15760);
   U10134 : AOI22_X1 port map( A1 => pipeline_data_to_RF_from_WB_13_port, A2 =>
                           n15605, B1 => pipeline_Alu_Out_Addr_to_mem_13_port, 
                           B2 => n17330, ZN => n15761);
   U10107 : AOI22_X1 port map( A1 => pipeline_stageF_PC_plus4_N26, A2 => n17108
                           , B1 => n17674, B2 => n13856, ZN => n15734);
   U10105 : AOI22_X1 port map( A1 => pipeline_stageD_target_Jump_temp_19_port, 
                           A2 => n17676, B1 => n17106, B2 => n15737, ZN => 
                           n15735);
   U10104 : AOI22_X1 port map( A1 => pipeline_data_to_RF_from_WB_19_port, A2 =>
                           n17333, B1 => pipeline_Alu_Out_Addr_to_mem_19_port, 
                           B2 => n17331, ZN => n15736);
   U10148 : AOI22_X1 port map( A1 => pipeline_stageF_PC_plus4_N7, A2 => n17108,
                           B1 => n17674, B2 => n13849, ZN => n15769);
   U10147 : AOI22_X1 port map( A1 => pipeline_stageD_target_Jump_temp_0_port, 
                           A2 => n17675, B1 => n17106, B2 => n15772, ZN => 
                           n15770);
   U10146 : AOI22_X1 port map( A1 => pipeline_data_to_RF_from_WB_0_port, A2 => 
                           n17333, B1 => pipeline_Alu_Out_Addr_to_mem_0_port, 
                           B2 => n15606, ZN => n15771);
   U10172 : AOI22_X1 port map( A1 => pipeline_stageF_PC_plus4_N12, A2 => n17108
                           , B1 => n17674, B2 => n13833, ZN => n15789);
   U10170 : AOI22_X1 port map( A1 => pipeline_stageD_target_Jump_temp_5_port, 
                           A2 => n15607, B1 => n17106, B2 => n15792, ZN => 
                           n15790);
   U10169 : AOI22_X1 port map( A1 => pipeline_data_to_RF_from_WB_5_port, A2 => 
                           n17333, B1 => pipeline_Alu_Out_Addr_to_mem_5_port, 
                           B2 => n17331, ZN => n15791);
   U10160 : AOI22_X1 port map( A1 => pipeline_stageF_PC_plus4_N14, A2 => n17108
                           , B1 => n17674, B2 => n13840, ZN => n15779);
   U10158 : AOI22_X1 port map( A1 => pipeline_stageD_target_Jump_temp_7_port, 
                           A2 => n17676, B1 => n17106, B2 => n15782, ZN => 
                           n15780);
   U10157 : AOI22_X1 port map( A1 => pipeline_data_to_RF_from_WB_7_port, A2 => 
                           n17333, B1 => pipeline_Alu_Out_Addr_to_mem_7_port, 
                           B2 => n17331, ZN => n15781);
   U10119 : AOI22_X1 port map( A1 => pipeline_stageF_PC_plus4_N24, A2 => n15610
                           , B1 => n17674, B2 => n13854, ZN => n15744);
   U10117 : AOI22_X1 port map( A1 => pipeline_stageD_target_Jump_temp_17_port, 
                           A2 => n15607, B1 => n17106, B2 => n15747, ZN => 
                           n15745);
   U10116 : AOI22_X1 port map( A1 => pipeline_data_to_RF_from_WB_17_port, A2 =>
                           n15605, B1 => pipeline_Alu_Out_Addr_to_mem_17_port, 
                           B2 => n15606, ZN => n15746);
   U10221 : AOI22_X1 port map( A1 => pipeline_stageF_PC_plus4_N8, A2 => n17108,
                           B1 => n17674, B2 => n13806, ZN => n15824);
   U10215 : AOI22_X1 port map( A1 => pipeline_stageD_target_Jump_temp_1_port, 
                           A2 => n17676, B1 => n17106, B2 => n15831, ZN => 
                           n15825);
   U10211 : AOI22_X1 port map( A1 => pipeline_data_to_RF_from_WB_1_port, A2 => 
                           n17332, B1 => pipeline_Alu_Out_Addr_to_mem_1_port, 
                           B2 => n17330, ZN => n15826);
   U10184 : AOI22_X1 port map( A1 => pipeline_stageF_PC_plus4_N18, A2 => n17108
                           , B1 => n17674, B2 => n13824, ZN => n15799);
   U10182 : AOI22_X1 port map( A1 => pipeline_stageD_target_Jump_temp_11_port, 
                           A2 => n17675, B1 => n17106, B2 => n15802, ZN => 
                           n15800);
   U10181 : AOI22_X1 port map( A1 => pipeline_data_to_RF_from_WB_11_port, A2 =>
                           n17332, B1 => pipeline_Alu_Out_Addr_to_mem_11_port, 
                           B2 => n17331, ZN => n15801);
   U10131 : AOI22_X1 port map( A1 => pipeline_stageF_PC_plus4_N21, A2 => n17108
                           , B1 => n17674, B2 => n13852, ZN => n15754);
   U10129 : AOI22_X1 port map( A1 => pipeline_stageD_target_Jump_temp_14_port, 
                           A2 => n17675, B1 => n17106, B2 => n15757, ZN => 
                           n15755);
   U10128 : AOI22_X1 port map( A1 => pipeline_data_to_RF_from_WB_14_port, A2 =>
                           n17333, B1 => pipeline_Alu_Out_Addr_to_mem_14_port, 
                           B2 => n17331, ZN => n15756);
   U10190 : AOI22_X1 port map( A1 => pipeline_stageF_PC_plus4_N16, A2 => n17108
                           , B1 => n17674, B2 => n13821, ZN => n15804);
   U10188 : AOI22_X1 port map( A1 => pipeline_stageD_target_Jump_temp_9_port, 
                           A2 => n15607, B1 => n15608, B2 => n15807, ZN => 
                           n15805);
   U10187 : AOI22_X1 port map( A1 => pipeline_data_to_RF_from_WB_9_port, A2 => 
                           n17332, B1 => pipeline_Alu_Out_Addr_to_mem_9_port, 
                           B2 => n17331, ZN => n15806);
   U9967 : AOI22_X1 port map( A1 => 
                           pipeline_stageD_offset_jump_sign_ext_24_port, A2 => 
                           n15600, B1 => n17672, B2 => InstrFetched_24_port, ZN
                           => n15644);
   U9935 : AOI22_X1 port map( A1 => n15600, A2 => 
                           pipeline_stageD_offset_to_jump_temp_7_port, B1 => 
                           n17672, B2 => InstrFetched_7_port, ZN => n15628);
   U9927 : AOI22_X1 port map( A1 => n15600, A2 => 
                           pipeline_stageD_offset_to_jump_temp_3_port, B1 => 
                           n17672, B2 => InstrFetched_3_port, ZN => n15624);
   U9911 : AOI22_X1 port map( A1 => n15600, A2 => 
                           pipeline_nextPC_IFID_DEC_16_port, B1 => n15601, B2 
                           => pipeline_stageF_PC_plus4_N23, ZN => n15612);
   U10180 : AOI22_X1 port map( A1 => n15600, A2 => 
                           pipeline_nextPC_IFID_DEC_6_port, B1 => n15601, B2 =>
                           pipeline_stageF_PC_plus4_N13, ZN => n15798);
   U10085 : AOI22_X1 port map( A1 => n15600, A2 => 
                           pipeline_nextPC_IFID_DEC_23_port, B1 => n15601, B2 
                           => pipeline_stageF_PC_plus4_N30, ZN => n15718);
   U9971 : AOI21_X1 port map( B1 => InstrFetched_26_port, B2 => n15646, A => 
                           n15648, ZN => n15647);
   U9970 : OAI21_X1 port map( B1 => n17409, B2 => n15646, A => n15647, ZN => 
                           n3962);
   U9979 : AOI21_X1 port map( B1 => InstrFetched_30_port, B2 => n15646, A => 
                           n15648, ZN => n15652);
   U9978 : OAI21_X1 port map( B1 => n17347, B2 => n15646, A => n15652, ZN => 
                           n3958);
   U9975 : AOI21_X1 port map( B1 => InstrFetched_28_port, B2 => n15646, A => 
                           n15648, ZN => n15650);
   U9974 : OAI21_X1 port map( B1 => n17348, B2 => n15646, A => n15650, ZN => 
                           n3960);
   U10987 : NAND2_X1 port map( A1 => n17701, A2 => 
                           pipeline_data_to_RF_from_WB_14_port, ZN => n15094);
   U9555 : OAI22_X1 port map( A1 => n17509, A2 => n17418, B1 => n17422, B2 => 
                           n15094, ZN => pipeline_EXMEM_stage_N53);
   U10965 : NAND2_X1 port map( A1 => n17702, A2 => 
                           pipeline_data_to_RF_from_WB_25_port, ZN => n15072);
   U9532 : OAI22_X1 port map( A1 => n17520, A2 => n17418, B1 => n17422, B2 => 
                           n15072, ZN => pipeline_EXMEM_stage_N64);
   U10979 : NAND2_X1 port map( A1 => n17702, A2 => 
                           pipeline_data_to_RF_from_WB_18_port, ZN => n15086);
   U9547 : OAI22_X1 port map( A1 => n17513, A2 => n17418, B1 => n17422, B2 => 
                           n15086, ZN => pipeline_EXMEM_stage_N57);
   U10973 : NAND2_X1 port map( A1 => n17702, A2 => 
                           pipeline_data_to_RF_from_WB_21_port, ZN => n15080);
   U9540 : OAI22_X1 port map( A1 => n17516, A2 => n17418, B1 => n17422, B2 => 
                           n15080, ZN => pipeline_EXMEM_stage_N60);
   U10955 : NAND2_X1 port map( A1 => n17703, A2 => 
                           pipeline_data_to_RF_from_WB_30_port, ZN => n15062);
   U9522 : OAI22_X1 port map( A1 => n17525, A2 => n17418, B1 => n17422, B2 => 
                           n15062, ZN => pipeline_EXMEM_stage_N69);
   U10999 : NAND2_X1 port map( A1 => n17704, A2 => 
                           pipeline_data_to_RF_from_WB_8_port, ZN => n15106);
   U9569 : OAI22_X1 port map( A1 => n17503, A2 => n17418, B1 => n17422, B2 => 
                           n15106, ZN => pipeline_EXMEM_stage_N47);
   U10953 : NAND2_X1 port map( A1 => n17703, A2 => 
                           pipeline_data_to_RF_from_WB_31_port, ZN => n14988);
   U9487 : OAI22_X1 port map( A1 => n17526, A2 => n17418, B1 => n17422, B2 => 
                           n14988, ZN => pipeline_EXMEM_stage_N70);
   U11005 : NAND2_X1 port map( A1 => n17704, A2 => 
                           pipeline_data_to_RF_from_WB_5_port, ZN => n15112);
   U9575 : OAI22_X1 port map( A1 => n17500, A2 => n17418, B1 => n17422, B2 => 
                           n15112, ZN => pipeline_EXMEM_stage_N44);
   U11001 : NAND2_X1 port map( A1 => n17704, A2 => 
                           pipeline_data_to_RF_from_WB_7_port, ZN => n15108);
   U9571 : OAI22_X1 port map( A1 => n17502, A2 => n17418, B1 => n17422, B2 => 
                           n15108, ZN => pipeline_EXMEM_stage_N46);
   U11011 : NAND2_X1 port map( A1 => n17704, A2 => 
                           pipeline_data_to_RF_from_WB_2_port, ZN => n15118);
   U9581 : OAI22_X1 port map( A1 => n17497, A2 => n17418, B1 => n17422, B2 => 
                           n15118, ZN => pipeline_EXMEM_stage_N41);
   U10975 : NAND2_X1 port map( A1 => n17701, A2 => 
                           pipeline_data_to_RF_from_WB_20_port, ZN => n15082);
   U9543 : OAI22_X1 port map( A1 => n17515, A2 => n17418, B1 => n17422, B2 => 
                           n15082, ZN => pipeline_EXMEM_stage_N59);
   U10991 : NAND2_X1 port map( A1 => n17704, A2 => 
                           pipeline_data_to_RF_from_WB_12_port, ZN => n15098);
   U9559 : OAI22_X1 port map( A1 => n17507, A2 => n17418, B1 => n17422, B2 => 
                           n15098, ZN => pipeline_EXMEM_stage_N51);
   U10985 : NAND2_X1 port map( A1 => n17702, A2 => 
                           pipeline_data_to_RF_from_WB_15_port, ZN => n15092);
   U9553 : OAI22_X1 port map( A1 => n17510, A2 => n17418, B1 => n17422, B2 => 
                           n15092, ZN => pipeline_EXMEM_stage_N54);
   U10995 : NAND2_X1 port map( A1 => n17704, A2 => 
                           pipeline_data_to_RF_from_WB_10_port, ZN => n15102);
   U9565 : OAI22_X1 port map( A1 => n17505, A2 => n17418, B1 => n17422, B2 => 
                           n15102, ZN => pipeline_EXMEM_stage_N49);
   U10997 : NAND2_X1 port map( A1 => n17704, A2 => 
                           pipeline_data_to_RF_from_WB_9_port, ZN => n15104);
   U9567 : OAI22_X1 port map( A1 => n17504, A2 => n17418, B1 => n17422, B2 => 
                           n15104, ZN => pipeline_EXMEM_stage_N48);
   U10981 : NAND2_X1 port map( A1 => n17701, A2 => 
                           pipeline_data_to_RF_from_WB_17_port, ZN => n15088);
   U9549 : OAI22_X1 port map( A1 => n17512, A2 => n17418, B1 => n17422, B2 => 
                           n15088, ZN => pipeline_EXMEM_stage_N56);
   U10969 : NAND2_X1 port map( A1 => n17701, A2 => 
                           pipeline_data_to_RF_from_WB_23_port, ZN => n15076);
   U9536 : OAI22_X1 port map( A1 => n17518, A2 => n17418, B1 => n17422, B2 => 
                           n15076, ZN => pipeline_EXMEM_stage_N62);
   U10983 : NAND2_X1 port map( A1 => n17702, A2 => 
                           pipeline_data_to_RF_from_WB_16_port, ZN => n15090);
   U9551 : OAI22_X1 port map( A1 => n17511, A2 => n17418, B1 => n17422, B2 => 
                           n15090, ZN => pipeline_EXMEM_stage_N55);
   U10977 : NAND2_X1 port map( A1 => n17701, A2 => 
                           pipeline_data_to_RF_from_WB_19_port, ZN => n15084);
   U9545 : OAI22_X1 port map( A1 => n17514, A2 => n17418, B1 => n17422, B2 => 
                           n15084, ZN => pipeline_EXMEM_stage_N58);
   U10963 : NAND2_X1 port map( A1 => n17702, A2 => 
                           pipeline_data_to_RF_from_WB_26_port, ZN => n15070);
   U9530 : OAI22_X1 port map( A1 => n17521, A2 => n17418, B1 => n17422, B2 => 
                           n15070, ZN => pipeline_EXMEM_stage_N65);
   U11007 : NAND2_X1 port map( A1 => n17704, A2 => 
                           pipeline_data_to_RF_from_WB_4_port, ZN => n15114);
   U9577 : OAI22_X1 port map( A1 => n17499, A2 => n17418, B1 => n17422, B2 => 
                           n15114, ZN => pipeline_EXMEM_stage_N43);
   U10989 : NAND2_X1 port map( A1 => n17704, A2 => 
                           pipeline_data_to_RF_from_WB_13_port, ZN => n15096);
   U9557 : OAI22_X1 port map( A1 => n17508, A2 => n17418, B1 => n17422, B2 => 
                           n15096, ZN => pipeline_EXMEM_stage_N52);
   U10959 : NAND2_X1 port map( A1 => n17703, A2 => 
                           pipeline_data_to_RF_from_WB_28_port, ZN => n15066);
   U9526 : OAI22_X1 port map( A1 => n17523, A2 => n17418, B1 => n17422, B2 => 
                           n15066, ZN => pipeline_EXMEM_stage_N67);
   U10967 : NAND2_X1 port map( A1 => n17701, A2 => 
                           pipeline_data_to_RF_from_WB_24_port, ZN => n15074);
   U9534 : OAI22_X1 port map( A1 => n17519, A2 => n17418, B1 => n17422, B2 => 
                           n15074, ZN => pipeline_EXMEM_stage_N63);
   U10971 : NAND2_X1 port map( A1 => n17701, A2 => 
                           pipeline_data_to_RF_from_WB_22_port, ZN => n15078);
   U9538 : OAI22_X1 port map( A1 => n17517, A2 => n17418, B1 => n17422, B2 => 
                           n15078, ZN => pipeline_EXMEM_stage_N61);
   U11003 : NAND2_X1 port map( A1 => n17704, A2 => 
                           pipeline_data_to_RF_from_WB_6_port, ZN => n15110);
   U9573 : OAI22_X1 port map( A1 => n17501, A2 => n17418, B1 => n17422, B2 => 
                           n15110, ZN => pipeline_EXMEM_stage_N45);
   U11013 : NAND2_X1 port map( A1 => n17704, A2 => 
                           pipeline_data_to_RF_from_WB_1_port, ZN => n15120);
   U9583 : OAI22_X1 port map( A1 => n17496, A2 => n17418, B1 => n17422, B2 => 
                           n15120, ZN => pipeline_EXMEM_stage_N40);
   U10957 : NAND2_X1 port map( A1 => n17703, A2 => 
                           pipeline_data_to_RF_from_WB_29_port, ZN => n15064);
   U9524 : OAI22_X1 port map( A1 => n17524, A2 => n17418, B1 => n17422, B2 => 
                           n15064, ZN => pipeline_EXMEM_stage_N68);
   U11015 : NAND2_X1 port map( A1 => n17704, A2 => 
                           pipeline_data_to_RF_from_WB_0_port, ZN => n15122);
   U9587 : OAI22_X1 port map( A1 => n17495, A2 => n17418, B1 => n17422, B2 => 
                           n15122, ZN => pipeline_EXMEM_stage_N39);
   U10961 : NAND2_X1 port map( A1 => n17703, A2 => 
                           pipeline_data_to_RF_from_WB_27_port, ZN => n15068);
   U9528 : OAI22_X1 port map( A1 => n17522, A2 => n17418, B1 => n17422, B2 => 
                           n15068, ZN => pipeline_EXMEM_stage_N66);
   U11009 : NAND2_X1 port map( A1 => n17703, A2 => 
                           pipeline_data_to_RF_from_WB_3_port, ZN => n15116);
   U9579 : OAI22_X1 port map( A1 => n17498, A2 => n17418, B1 => n17422, B2 => 
                           n15116, ZN => pipeline_EXMEM_stage_N42);
   U10993 : NAND2_X1 port map( A1 => n17704, A2 => 
                           pipeline_data_to_RF_from_WB_11_port, ZN => n15100);
   U9561 : OAI22_X1 port map( A1 => n17506, A2 => n17418, B1 => n17422, B2 => 
                           n15100, ZN => pipeline_EXMEM_stage_N50);
   U8678 : NOR2_X1 port map( A1 => n17431, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N181);
   U8989 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_31_18_port,
                           A2 => n17154, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_18_port, B2 => 
                           n17683, ZN => n14508);
   U8988 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_29_18_port,
                           A2 => n17684, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_18_port, B2 => 
                           n17685, ZN => n14509);
   U9375 : NAND2_X1 port map( A1 => n17408, A2 => n17329, ZN => n14860);
   U8987 : AOI222_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_4_18_port,
                           A2 => n17686, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_18_port, B2 => 
                           n17153, C1 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_18_port, C2 => 
                           n17687, ZN => n14510);
   U8986 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_27_18_port,
                           A2 => n17688, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_18_port, B2 => 
                           n17689, ZN => n14504);
   U8985 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_23_18_port,
                           A2 => n17690, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_18_port, B2 => 
                           n17691, ZN => n14505);
   U8984 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_21_18_port,
                           A2 => n17692, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_18_port, B2 => 
                           n17693, ZN => n14506);
   U8983 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_19_18_port,
                           A2 => n17694, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_18_port, B2 => 
                           n17695, ZN => n14507);
   U8982 : NAND4_X1 port map( A1 => n14504, A2 => n14505, A3 => n14506, A4 => 
                           n14507, ZN => n14493);
   U8981 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_17_18_port,
                           A2 => n17696, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_18_port, B2 => 
                           n17697, ZN => n14500);
   U9353 : NOR2_X1 port map( A1 => n14865, A2 => n14867, ZN => n14226);
   U8980 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_12_18_port,
                           A2 => n17698, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_18_port, B2 => 
                           n14226, ZN => n14501);
   U8979 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_8_18_port, 
                           A2 => n14223, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_18_port, B2 => 
                           n17152, ZN => n14502);
   U9348 : NOR2_X1 port map( A1 => n14860, A2 => n14867, ZN => n14221);
   U8978 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_9_18_port, 
                           A2 => n14221, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_18_port, B2 => 
                           n17699, ZN => n14503);
   U8977 : NAND4_X1 port map( A1 => n14500, A2 => n14501, A3 => n14502, A4 => 
                           n14503, ZN => n14494);
   U8976 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_11_18_port,
                           A2 => n17151, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_18_port, B2 => 
                           n14216, ZN => n14496);
   U8975 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_14_18_port,
                           A2 => n17700, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_18_port, B2 => 
                           n14214, ZN => n14497);
   U8974 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_2_18_port, 
                           A2 => n17367, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_18_port, B2 => 
                           n14212, ZN => n14498);
   U8973 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_6_18_port, 
                           A2 => n17368, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_18_port, B2 => 
                           n14210, ZN => n14499);
   U8972 : NAND4_X1 port map( A1 => n14496, A2 => n14497, A3 => n14498, A4 => 
                           n14499, ZN => n14495);
   U8971 : NOR4_X1 port map( A1 => n14492, A2 => n14493, A3 => n14494, A4 => 
                           n14495, ZN => n14491);
   U8970 : NOR2_X1 port map( A1 => n14491, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N152);
   U9229 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_31_6_port, 
                           A2 => n17154, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_6_port, B2 => 
                           n17683, ZN => n14748);
   U9228 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_29_6_port, 
                           A2 => n17684, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_6_port, B2 => 
                           n17685, ZN => n14749);
   U9227 : AOI222_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_4_6_port, 
                           A2 => n17686, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_6_port, B2 => 
                           n17153, C1 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_6_port, C2 => 
                           n17687, ZN => n14750);
   U9226 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_27_6_port, 
                           A2 => n17688, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_6_port, B2 => 
                           n17689, ZN => n14744);
   U9225 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_23_6_port, 
                           A2 => n17690, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_6_port, B2 => 
                           n17691, ZN => n14745);
   U9224 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_21_6_port, 
                           A2 => n17692, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_6_port, B2 => 
                           n17693, ZN => n14746);
   U9223 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_19_6_port, 
                           A2 => n17694, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_6_port, B2 => 
                           n17695, ZN => n14747);
   U9222 : NAND4_X1 port map( A1 => n14744, A2 => n14745, A3 => n14746, A4 => 
                           n14747, ZN => n14733);
   U9221 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_17_6_port, 
                           A2 => n17696, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_6_port, B2 => 
                           n17697, ZN => n14740);
   U9220 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_12_6_port, 
                           A2 => n17698, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_6_port, B2 => 
                           n17358, ZN => n14741);
   U9219 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_8_6_port, 
                           A2 => n17417, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_6_port, B2 => 
                           n17152, ZN => n14742);
   U9218 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_9_6_port, 
                           A2 => n17352, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_6_port, B2 => 
                           n17699, ZN => n14743);
   U9217 : NAND4_X1 port map( A1 => n14740, A2 => n14741, A3 => n14742, A4 => 
                           n14743, ZN => n14734);
   U9216 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_11_6_port, 
                           A2 => n17151, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_6_port, B2 => 
                           n17413, ZN => n14736);
   U9215 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_14_6_port, 
                           A2 => n17700, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_6_port, B2 => 
                           n17414, ZN => n14737);
   U9214 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_2_6_port, 
                           A2 => n17355, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_6_port, B2 => 
                           n17415, ZN => n14738);
   U9213 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_6_6_port, 
                           A2 => n17356, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_6_port, B2 => 
                           n17416, ZN => n14739);
   U9212 : NAND4_X1 port map( A1 => n14736, A2 => n14737, A3 => n14738, A4 => 
                           n14739, ZN => n14735);
   U9211 : NOR4_X1 port map( A1 => n14732, A2 => n14733, A3 => n14734, A4 => 
                           n14735, ZN => n14731);
   U9210 : NOR2_X1 port map( A1 => n14731, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N140);
   U9169 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_31_9_port, 
                           A2 => n17154, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_9_port, B2 => 
                           n17683, ZN => n14688);
   U9168 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_29_9_port, 
                           A2 => n17684, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_9_port, B2 => 
                           n17685, ZN => n14689);
   U9167 : AOI222_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_4_9_port, 
                           A2 => n17686, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_9_port, B2 => 
                           n17153, C1 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_9_port, C2 => 
                           n14246, ZN => n14690);
   U9166 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_27_9_port, 
                           A2 => n17688, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_9_port, B2 => 
                           n17689, ZN => n14684);
   U9165 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_23_9_port, 
                           A2 => n17690, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_9_port, B2 => 
                           n17691, ZN => n14685);
   U9164 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_21_9_port, 
                           A2 => n17692, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_9_port, B2 => 
                           n17693, ZN => n14686);
   U9163 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_19_9_port, 
                           A2 => n17694, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_9_port, B2 => 
                           n17695, ZN => n14687);
   U9162 : NAND4_X1 port map( A1 => n14684, A2 => n14685, A3 => n14686, A4 => 
                           n14687, ZN => n14673);
   U9161 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_17_9_port, 
                           A2 => n17696, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_9_port, B2 => 
                           n17697, ZN => n14680);
   U9160 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_12_9_port, 
                           A2 => n17698, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_9_port, B2 => 
                           n17358, ZN => n14681);
   U9159 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_8_9_port, 
                           A2 => n14223, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_9_port, B2 => 
                           n17152, ZN => n14682);
   U9158 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_9_9_port, 
                           A2 => n17352, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_9_port, B2 => 
                           n17699, ZN => n14683);
   U9157 : NAND4_X1 port map( A1 => n14680, A2 => n14681, A3 => n14682, A4 => 
                           n14683, ZN => n14674);
   U9156 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_11_9_port, 
                           A2 => n17151, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_9_port, B2 => 
                           n14216, ZN => n14676);
   U9155 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_14_9_port, 
                           A2 => n17700, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_9_port, B2 => 
                           n14214, ZN => n14677);
   U9154 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_2_9_port, 
                           A2 => n17355, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_9_port, B2 => 
                           n14212, ZN => n14678);
   U9153 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_6_9_port, 
                           A2 => n17356, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_9_port, B2 => 
                           n14210, ZN => n14679);
   U9152 : NAND4_X1 port map( A1 => n14676, A2 => n14677, A3 => n14678, A4 => 
                           n14679, ZN => n14675);
   U9151 : NOR4_X1 port map( A1 => n14672, A2 => n14673, A3 => n14674, A4 => 
                           n14675, ZN => n14671);
   U9150 : NOR2_X1 port map( A1 => n14671, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N143);
   U8809 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_31_27_port,
                           A2 => n14249, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_27_port, B2 => 
                           n14250, ZN => n14328);
   U8808 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_29_27_port,
                           A2 => n14247, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_27_port, B2 => 
                           n14248, ZN => n14329);
   U8807 : AOI222_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_4_27_port,
                           A2 => n14244, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_27_port, B2 => 
                           n14245, C1 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_27_port, C2 => 
                           n17687, ZN => n14330);
   U8806 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_27_27_port,
                           A2 => n14239, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_27_port, B2 => 
                           n14240, ZN => n14324);
   U8805 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_23_27_port,
                           A2 => n14237, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_27_port, B2 => 
                           n14238, ZN => n14325);
   U8804 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_21_27_port,
                           A2 => n14235, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_27_port, B2 => 
                           n14236, ZN => n14326);
   U8803 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_19_27_port,
                           A2 => n14233, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_27_port, B2 => 
                           n14234, ZN => n14327);
   U8802 : NAND4_X1 port map( A1 => n14324, A2 => n14325, A3 => n14326, A4 => 
                           n14327, ZN => n14313);
   U8801 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_17_27_port,
                           A2 => n14227, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_27_port, B2 => 
                           n14228, ZN => n14320);
   U8800 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_12_27_port,
                           A2 => n14225, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_27_port, B2 => 
                           n17357, ZN => n14321);
   U8799 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_8_27_port, 
                           A2 => n17417, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_27_port, B2 => 
                           n17152, ZN => n14322);
   U8798 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_9_27_port, 
                           A2 => n17351, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_27_port, B2 => 
                           n14222, ZN => n14323);
   U8797 : NAND4_X1 port map( A1 => n14320, A2 => n14321, A3 => n14322, A4 => 
                           n14323, ZN => n14314);
   U8796 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_11_27_port,
                           A2 => n17151, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_27_port, B2 => 
                           n17413, ZN => n14316);
   U8795 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_14_27_port,
                           A2 => n17700, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_27_port, B2 => 
                           n17414, ZN => n14317);
   U8794 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_2_27_port, 
                           A2 => n17353, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_27_port, B2 => 
                           n17415, ZN => n14318);
   U8793 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_6_27_port, 
                           A2 => n17354, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_27_port, B2 => 
                           n17416, ZN => n14319);
   U8792 : NAND4_X1 port map( A1 => n14316, A2 => n14317, A3 => n14318, A4 => 
                           n14319, ZN => n14315);
   U8791 : NOR4_X1 port map( A1 => n14312, A2 => n14313, A3 => n14314, A4 => 
                           n14315, ZN => n14311);
   U8790 : NOR2_X1 port map( A1 => n14311, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N161);
   U8969 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_31_19_port,
                           A2 => n17154, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_19_port, B2 => 
                           n17683, ZN => n14488);
   U8968 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_29_19_port,
                           A2 => n17684, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_19_port, B2 => 
                           n17685, ZN => n14489);
   U8967 : AOI222_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_4_19_port,
                           A2 => n17686, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_19_port, B2 => 
                           n17153, C1 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_19_port, C2 => 
                           n17687, ZN => n14490);
   U8966 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_27_19_port,
                           A2 => n17688, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_19_port, B2 => 
                           n17689, ZN => n14484);
   U8965 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_23_19_port,
                           A2 => n17690, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_19_port, B2 => 
                           n17691, ZN => n14485);
   U8964 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_21_19_port,
                           A2 => n17692, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_19_port, B2 => 
                           n17693, ZN => n14486);
   U8963 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_19_19_port,
                           A2 => n17694, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_19_port, B2 => 
                           n17695, ZN => n14487);
   U8962 : NAND4_X1 port map( A1 => n14484, A2 => n14485, A3 => n14486, A4 => 
                           n14487, ZN => n14473);
   U8961 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_17_19_port,
                           A2 => n17696, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_19_port, B2 => 
                           n17697, ZN => n14480);
   U8960 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_12_19_port,
                           A2 => n17698, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_19_port, B2 => 
                           n14226, ZN => n14481);
   U8959 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_8_19_port, 
                           A2 => n14223, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_19_port, B2 => 
                           n17152, ZN => n14482);
   U8958 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_9_19_port, 
                           A2 => n14221, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_19_port, B2 => 
                           n17699, ZN => n14483);
   U8957 : NAND4_X1 port map( A1 => n14480, A2 => n14481, A3 => n14482, A4 => 
                           n14483, ZN => n14474);
   U8956 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_11_19_port,
                           A2 => n17151, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_19_port, B2 => 
                           n14216, ZN => n14476);
   U8955 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_14_19_port,
                           A2 => n17700, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_19_port, B2 => 
                           n14214, ZN => n14477);
   U8954 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_2_19_port, 
                           A2 => n17367, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_19_port, B2 => 
                           n14212, ZN => n14478);
   U8953 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_6_19_port, 
                           A2 => n17368, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_19_port, B2 => 
                           n14210, ZN => n14479);
   U8952 : NAND4_X1 port map( A1 => n14476, A2 => n14477, A3 => n14478, A4 => 
                           n14479, ZN => n14475);
   U8951 : NOR4_X1 port map( A1 => n14472, A2 => n14473, A3 => n14474, A4 => 
                           n14475, ZN => n14471);
   U8950 : NOR2_X1 port map( A1 => n14471, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N153);
   U9049 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_31_15_port,
                           A2 => n17154, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_15_port, B2 => 
                           n17683, ZN => n14568);
   U9048 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_29_15_port,
                           A2 => n17684, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_15_port, B2 => 
                           n17685, ZN => n14569);
   U9047 : AOI222_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_4_15_port,
                           A2 => n17686, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_15_port, B2 => 
                           n17153, C1 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_15_port, C2 => 
                           n17687, ZN => n14570);
   U9046 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_27_15_port,
                           A2 => n17688, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_15_port, B2 => 
                           n17689, ZN => n14564);
   U9045 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_23_15_port,
                           A2 => n17690, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_15_port, B2 => 
                           n17691, ZN => n14565);
   U9044 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_21_15_port,
                           A2 => n17692, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_15_port, B2 => 
                           n17693, ZN => n14566);
   U9043 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_19_15_port,
                           A2 => n17694, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_15_port, B2 => 
                           n17695, ZN => n14567);
   U9042 : NAND4_X1 port map( A1 => n14564, A2 => n14565, A3 => n14566, A4 => 
                           n14567, ZN => n14553);
   U9041 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_17_15_port,
                           A2 => n17696, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_15_port, B2 => 
                           n17697, ZN => n14560);
   U9040 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_12_15_port,
                           A2 => n17698, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_15_port, B2 => 
                           n17358, ZN => n14561);
   U9039 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_8_15_port, 
                           A2 => n14223, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_15_port, B2 => 
                           n17152, ZN => n14562);
   U9038 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_9_15_port, 
                           A2 => n17352, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_15_port, B2 => 
                           n17699, ZN => n14563);
   U9037 : NAND4_X1 port map( A1 => n14560, A2 => n14561, A3 => n14562, A4 => 
                           n14563, ZN => n14554);
   U9036 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_11_15_port,
                           A2 => n17151, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_15_port, B2 => 
                           n14216, ZN => n14556);
   U9035 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_14_15_port,
                           A2 => n17700, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_15_port, B2 => 
                           n14214, ZN => n14557);
   U9034 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_2_15_port, 
                           A2 => n17355, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_15_port, B2 => 
                           n14212, ZN => n14558);
   U9033 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_6_15_port, 
                           A2 => n17356, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_15_port, B2 => 
                           n14210, ZN => n14559);
   U9032 : NAND4_X1 port map( A1 => n14556, A2 => n14557, A3 => n14558, A4 => 
                           n14559, ZN => n14555);
   U9031 : NOR4_X1 port map( A1 => n14552, A2 => n14553, A3 => n14554, A4 => 
                           n14555, ZN => n14551);
   U9030 : NOR2_X1 port map( A1 => n14551, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N149);
   U9009 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_31_17_port,
                           A2 => n17154, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_17_port, B2 => 
                           n17683, ZN => n14528);
   U9008 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_29_17_port,
                           A2 => n17684, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_17_port, B2 => 
                           n17685, ZN => n14529);
   U9007 : AOI222_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_4_17_port,
                           A2 => n17686, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_17_port, B2 => 
                           n17153, C1 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_17_port, C2 => 
                           n17687, ZN => n14530);
   U9006 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_27_17_port,
                           A2 => n17688, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_17_port, B2 => 
                           n17689, ZN => n14524);
   U9005 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_23_17_port,
                           A2 => n17690, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_17_port, B2 => 
                           n17691, ZN => n14525);
   U9004 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_21_17_port,
                           A2 => n17692, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_17_port, B2 => 
                           n17693, ZN => n14526);
   U9003 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_19_17_port,
                           A2 => n17694, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_17_port, B2 => 
                           n17695, ZN => n14527);
   U9002 : NAND4_X1 port map( A1 => n14524, A2 => n14525, A3 => n14526, A4 => 
                           n14527, ZN => n14513);
   U9001 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_17_17_port,
                           A2 => n17696, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_17_port, B2 => 
                           n17697, ZN => n14520);
   U9000 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_12_17_port,
                           A2 => n17698, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_17_port, B2 => 
                           n14226, ZN => n14521);
   U8999 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_8_17_port, 
                           A2 => n14223, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_17_port, B2 => 
                           n17152, ZN => n14522);
   U8998 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_9_17_port, 
                           A2 => n14221, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_17_port, B2 => 
                           n17699, ZN => n14523);
   U8997 : NAND4_X1 port map( A1 => n14520, A2 => n14521, A3 => n14522, A4 => 
                           n14523, ZN => n14514);
   U8996 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_11_17_port,
                           A2 => n17151, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_17_port, B2 => 
                           n14216, ZN => n14516);
   U8995 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_14_17_port,
                           A2 => n17700, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_17_port, B2 => 
                           n14214, ZN => n14517);
   U8994 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_2_17_port, 
                           A2 => n17367, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_17_port, B2 => 
                           n14212, ZN => n14518);
   U8993 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_6_17_port, 
                           A2 => n17368, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_17_port, B2 => 
                           n14210, ZN => n14519);
   U8992 : NAND4_X1 port map( A1 => n14516, A2 => n14517, A3 => n14518, A4 => 
                           n14519, ZN => n14515);
   U8991 : NOR4_X1 port map( A1 => n14512, A2 => n14513, A3 => n14514, A4 => 
                           n14515, ZN => n14511);
   U8990 : NOR2_X1 port map( A1 => n14511, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N151);
   U9385 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_31_0_port, 
                           A2 => n14249, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_0_port, B2 => 
                           n14250, ZN => n14880);
   U9380 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_29_0_port, 
                           A2 => n14247, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_0_port, B2 => 
                           n14248, ZN => n14881);
   U9372 : AOI222_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_4_0_port, 
                           A2 => n14244, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_0_port, B2 => 
                           n17153, C1 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_0_port, C2 => 
                           n17687, ZN => n14882);
   U9368 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_27_0_port, 
                           A2 => n14239, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_0_port, B2 => 
                           n14240, ZN => n14874);
   U9365 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_23_0_port, 
                           A2 => n14237, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_0_port, B2 => 
                           n14238, ZN => n14875);
   U9362 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_21_0_port, 
                           A2 => n14235, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_0_port, B2 => 
                           n14236, ZN => n14876);
   U9359 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_19_0_port, 
                           A2 => n14233, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_0_port, B2 => 
                           n14234, ZN => n14877);
   U9358 : NAND4_X1 port map( A1 => n14874, A2 => n14875, A3 => n14876, A4 => 
                           n14877, ZN => n14853);
   U9355 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_17_0_port, 
                           A2 => n14227, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_0_port, B2 => 
                           n14228, ZN => n14868);
   U9352 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_12_0_port, 
                           A2 => n14225, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_0_port, B2 => 
                           n17357, ZN => n14869);
   U9349 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_8_0_port, 
                           A2 => n17417, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_0_port, B2 => 
                           n17152, ZN => n14870);
   U9346 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_9_0_port, 
                           A2 => n17351, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_0_port, B2 => 
                           n14222, ZN => n14871);
   U9345 : NAND4_X1 port map( A1 => n14868, A2 => n14869, A3 => n14870, A4 => 
                           n14871, ZN => n14854);
   U9342 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_11_0_port, 
                           A2 => n17151, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_0_port, B2 => 
                           n17413, ZN => n14856);
   U9339 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_14_0_port, 
                           A2 => n17700, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_0_port, B2 => 
                           n17414, ZN => n14857);
   U9336 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_2_0_port, 
                           A2 => n17353, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_0_port, B2 => 
                           n17415, ZN => n14858);
   U9333 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_6_0_port, 
                           A2 => n17354, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_0_port, B2 => 
                           n17416, ZN => n14859);
   U9332 : NAND4_X1 port map( A1 => n14856, A2 => n14857, A3 => n14858, A4 => 
                           n14859, ZN => n14855);
   U9331 : NOR4_X1 port map( A1 => n14852, A2 => n14853, A3 => n14854, A4 => 
                           n14855, ZN => n14851);
   U9330 : NOR2_X1 port map( A1 => n14851, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N134);
   U9269 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_31_4_port, 
                           A2 => n17154, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_4_port, B2 => 
                           n17683, ZN => n14788);
   U9268 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_29_4_port, 
                           A2 => n17684, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_4_port, B2 => 
                           n17685, ZN => n14789);
   U9267 : AOI222_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_4_4_port, 
                           A2 => n17686, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_4_port, B2 => 
                           n17153, C1 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_4_port, C2 => 
                           n14246, ZN => n14790);
   U9266 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_27_4_port, 
                           A2 => n17688, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_4_port, B2 => 
                           n17689, ZN => n14784);
   U9265 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_23_4_port, 
                           A2 => n17690, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_4_port, B2 => 
                           n17691, ZN => n14785);
   U9264 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_21_4_port, 
                           A2 => n17692, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_4_port, B2 => 
                           n17693, ZN => n14786);
   U9263 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_19_4_port, 
                           A2 => n17694, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_4_port, B2 => 
                           n17695, ZN => n14787);
   U9262 : NAND4_X1 port map( A1 => n14784, A2 => n14785, A3 => n14786, A4 => 
                           n14787, ZN => n14773);
   U9261 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_17_4_port, 
                           A2 => n17696, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_4_port, B2 => 
                           n17697, ZN => n14780);
   U9260 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_12_4_port, 
                           A2 => n17698, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_4_port, B2 => 
                           n17357, ZN => n14781);
   U9259 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_8_4_port, 
                           A2 => n17417, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_4_port, B2 => 
                           n17152, ZN => n14782);
   U9258 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_9_4_port, 
                           A2 => n17351, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_4_port, B2 => 
                           n17699, ZN => n14783);
   U9257 : NAND4_X1 port map( A1 => n14780, A2 => n14781, A3 => n14782, A4 => 
                           n14783, ZN => n14774);
   U9256 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_11_4_port, 
                           A2 => n14215, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_4_port, B2 => 
                           n17413, ZN => n14776);
   U9255 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_14_4_port, 
                           A2 => n17700, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_4_port, B2 => 
                           n17414, ZN => n14777);
   U9254 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_2_4_port, 
                           A2 => n17353, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_4_port, B2 => 
                           n17415, ZN => n14778);
   U9253 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_6_4_port, 
                           A2 => n17354, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_4_port, B2 => 
                           n17416, ZN => n14779);
   U9252 : NAND4_X1 port map( A1 => n14776, A2 => n14777, A3 => n14778, A4 => 
                           n14779, ZN => n14775);
   U9251 : NOR4_X1 port map( A1 => n14772, A2 => n14773, A3 => n14774, A4 => 
                           n14775, ZN => n14771);
   U9250 : NOR2_X1 port map( A1 => n14771, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N138);
   U8909 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_31_22_port,
                           A2 => n17154, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_22_port, B2 => 
                           n17683, ZN => n14428);
   U8908 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_29_22_port,
                           A2 => n17684, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_22_port, B2 => 
                           n17685, ZN => n14429);
   U8907 : AOI222_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_4_22_port,
                           A2 => n17686, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_22_port, B2 => 
                           n14245, C1 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_22_port, C2 => 
                           n14246, ZN => n14430);
   U8906 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_27_22_port,
                           A2 => n14239, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_22_port, B2 => 
                           n17689, ZN => n14424);
   U8905 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_23_22_port,
                           A2 => n17690, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_22_port, B2 => 
                           n17691, ZN => n14425);
   U8904 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_21_22_port,
                           A2 => n14235, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_22_port, B2 => 
                           n17693, ZN => n14426);
   U8903 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_19_22_port,
                           A2 => n17694, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_22_port, B2 => 
                           n17695, ZN => n14427);
   U8902 : NAND4_X1 port map( A1 => n14424, A2 => n14425, A3 => n14426, A4 => 
                           n14427, ZN => n14413);
   U8901 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_17_22_port,
                           A2 => n14227, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_22_port, B2 => 
                           n17697, ZN => n14420);
   U8900 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_12_22_port,
                           A2 => n17698, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_22_port, B2 => 
                           n17357, ZN => n14421);
   U8899 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_8_22_port, 
                           A2 => n17417, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_22_port, B2 => 
                           n17152, ZN => n14422);
   U8898 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_9_22_port, 
                           A2 => n17351, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_22_port, B2 => 
                           n17699, ZN => n14423);
   U8897 : NAND4_X1 port map( A1 => n14420, A2 => n14421, A3 => n14422, A4 => 
                           n14423, ZN => n14414);
   U8896 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_11_22_port,
                           A2 => n14215, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_22_port, B2 => 
                           n17413, ZN => n14416);
   U8895 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_14_22_port,
                           A2 => n14213, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_22_port, B2 => 
                           n17414, ZN => n14417);
   U8894 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_2_22_port, 
                           A2 => n17353, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_22_port, B2 => 
                           n17415, ZN => n14418);
   U8893 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_6_22_port, 
                           A2 => n17354, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_22_port, B2 => 
                           n17416, ZN => n14419);
   U8892 : NAND4_X1 port map( A1 => n14416, A2 => n14417, A3 => n14418, A4 => 
                           n14419, ZN => n14415);
   U8891 : NOR4_X1 port map( A1 => n14412, A2 => n14413, A3 => n14414, A4 => 
                           n14415, ZN => n14411);
   U8890 : NOR2_X1 port map( A1 => n14411, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N156);
   U9249 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_31_5_port, 
                           A2 => n17154, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_5_port, B2 => 
                           n17683, ZN => n14768);
   U9248 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_29_5_port, 
                           A2 => n17684, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_5_port, B2 => 
                           n17685, ZN => n14769);
   U9247 : AOI222_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_4_5_port, 
                           A2 => n17686, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_5_port, B2 => 
                           n17153, C1 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_5_port, C2 => 
                           n17687, ZN => n14770);
   U9246 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_27_5_port, 
                           A2 => n17688, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_5_port, B2 => 
                           n17689, ZN => n14764);
   U9245 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_23_5_port, 
                           A2 => n17690, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_5_port, B2 => 
                           n17691, ZN => n14765);
   U9244 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_21_5_port, 
                           A2 => n17692, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_5_port, B2 => 
                           n17693, ZN => n14766);
   U9243 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_19_5_port, 
                           A2 => n17694, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_5_port, B2 => 
                           n17695, ZN => n14767);
   U9242 : NAND4_X1 port map( A1 => n14764, A2 => n14765, A3 => n14766, A4 => 
                           n14767, ZN => n14753);
   U9241 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_17_5_port, 
                           A2 => n17696, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_5_port, B2 => 
                           n17697, ZN => n14760);
   U9240 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_12_5_port, 
                           A2 => n17698, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_5_port, B2 => 
                           n17357, ZN => n14761);
   U9239 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_8_5_port, 
                           A2 => n17417, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_5_port, B2 => 
                           n17152, ZN => n14762);
   U9238 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_9_5_port, 
                           A2 => n17351, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_5_port, B2 => 
                           n17699, ZN => n14763);
   U9237 : NAND4_X1 port map( A1 => n14760, A2 => n14761, A3 => n14762, A4 => 
                           n14763, ZN => n14754);
   U9236 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_11_5_port, 
                           A2 => n14215, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_5_port, B2 => 
                           n17413, ZN => n14756);
   U9235 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_14_5_port, 
                           A2 => n17700, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_5_port, B2 => 
                           n17414, ZN => n14757);
   U9234 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_2_5_port, 
                           A2 => n17353, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_5_port, B2 => 
                           n17415, ZN => n14758);
   U9233 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_6_5_port, 
                           A2 => n17354, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_5_port, B2 => 
                           n17416, ZN => n14759);
   U9232 : NAND4_X1 port map( A1 => n14756, A2 => n14757, A3 => n14758, A4 => 
                           n14759, ZN => n14755);
   U9231 : NOR4_X1 port map( A1 => n14752, A2 => n14753, A3 => n14754, A4 => 
                           n14755, ZN => n14751);
   U9230 : NOR2_X1 port map( A1 => n14751, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N139);
   U8889 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_31_23_port,
                           A2 => n14249, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_23_port, B2 => 
                           n17683, ZN => n14408);
   U8888 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_29_23_port,
                           A2 => n17684, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_23_port, B2 => 
                           n17685, ZN => n14409);
   U8887 : AOI222_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_4_23_port,
                           A2 => n17686, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_23_port, B2 => 
                           n14245, C1 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_23_port, C2 => 
                           n17687, ZN => n14410);
   U8886 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_27_23_port,
                           A2 => n14239, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_23_port, B2 => 
                           n17689, ZN => n14404);
   U8885 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_23_23_port,
                           A2 => n14237, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_23_port, B2 => 
                           n17691, ZN => n14405);
   U8884 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_21_23_port,
                           A2 => n17692, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_23_port, B2 => 
                           n17693, ZN => n14406);
   U8883 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_19_23_port,
                           A2 => n17694, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_23_port, B2 => 
                           n17695, ZN => n14407);
   U8882 : NAND4_X1 port map( A1 => n14404, A2 => n14405, A3 => n14406, A4 => 
                           n14407, ZN => n14393);
   U8881 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_17_23_port,
                           A2 => n14227, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_23_port, B2 => 
                           n17697, ZN => n14400);
   U8880 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_12_23_port,
                           A2 => n17698, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_23_port, B2 => 
                           n17357, ZN => n14401);
   U8879 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_8_23_port, 
                           A2 => n17417, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_23_port, B2 => 
                           n17152, ZN => n14402);
   U8878 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_9_23_port, 
                           A2 => n17351, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_23_port, B2 => 
                           n17699, ZN => n14403);
   U8877 : NAND4_X1 port map( A1 => n14400, A2 => n14401, A3 => n14402, A4 => 
                           n14403, ZN => n14394);
   U8876 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_11_23_port,
                           A2 => n14215, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_23_port, B2 => 
                           n17413, ZN => n14396);
   U8875 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_14_23_port,
                           A2 => n14213, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_23_port, B2 => 
                           n17414, ZN => n14397);
   U8874 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_2_23_port, 
                           A2 => n17353, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_23_port, B2 => 
                           n17415, ZN => n14398);
   U8873 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_6_23_port, 
                           A2 => n17354, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_23_port, B2 => 
                           n17416, ZN => n14399);
   U8872 : NAND4_X1 port map( A1 => n14396, A2 => n14397, A3 => n14398, A4 => 
                           n14399, ZN => n14395);
   U8871 : NOR4_X1 port map( A1 => n14392, A2 => n14393, A3 => n14394, A4 => 
                           n14395, ZN => n14391);
   U8870 : NOR2_X1 port map( A1 => n14391, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N157);
   U9089 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_31_13_port,
                           A2 => n17154, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_13_port, B2 => 
                           n17683, ZN => n14608);
   U9088 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_29_13_port,
                           A2 => n17684, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_13_port, B2 => 
                           n17685, ZN => n14609);
   U9087 : AOI222_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_4_13_port,
                           A2 => n17686, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_13_port, B2 => 
                           n17153, C1 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_13_port, C2 => 
                           n17687, ZN => n14610);
   U9086 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_27_13_port,
                           A2 => n17688, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_13_port, B2 => 
                           n17689, ZN => n14604);
   U9085 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_23_13_port,
                           A2 => n17690, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_13_port, B2 => 
                           n17691, ZN => n14605);
   U9084 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_21_13_port,
                           A2 => n17692, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_13_port, B2 => 
                           n17693, ZN => n14606);
   U9083 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_19_13_port,
                           A2 => n17694, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_13_port, B2 => 
                           n17695, ZN => n14607);
   U9082 : NAND4_X1 port map( A1 => n14604, A2 => n14605, A3 => n14606, A4 => 
                           n14607, ZN => n14593);
   U9081 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_17_13_port,
                           A2 => n17696, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_13_port, B2 => 
                           n17697, ZN => n14600);
   U9080 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_12_13_port,
                           A2 => n17698, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_13_port, B2 => 
                           n14226, ZN => n14601);
   U9079 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_8_13_port, 
                           A2 => n14223, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_13_port, B2 => 
                           n17152, ZN => n14602);
   U9078 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_9_13_port, 
                           A2 => n14221, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_13_port, B2 => 
                           n17699, ZN => n14603);
   U9077 : NAND4_X1 port map( A1 => n14600, A2 => n14601, A3 => n14602, A4 => 
                           n14603, ZN => n14594);
   U9076 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_11_13_port,
                           A2 => n17151, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_13_port, B2 => 
                           n14216, ZN => n14596);
   U9075 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_14_13_port,
                           A2 => n17700, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_13_port, B2 => 
                           n14214, ZN => n14597);
   U9074 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_2_13_port, 
                           A2 => n17367, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_13_port, B2 => 
                           n14212, ZN => n14598);
   U9073 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_6_13_port, 
                           A2 => n17368, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_13_port, B2 => 
                           n14210, ZN => n14599);
   U9072 : NAND4_X1 port map( A1 => n14596, A2 => n14597, A3 => n14598, A4 => 
                           n14599, ZN => n14595);
   U9071 : NOR4_X1 port map( A1 => n14592, A2 => n14593, A3 => n14594, A4 => 
                           n14595, ZN => n14591);
   U9070 : NOR2_X1 port map( A1 => n14591, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N147);
   U9069 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_31_14_port,
                           A2 => n17154, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_14_port, B2 => 
                           n17683, ZN => n14588);
   U9068 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_29_14_port,
                           A2 => n17684, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_14_port, B2 => 
                           n17685, ZN => n14589);
   U9067 : AOI222_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_4_14_port,
                           A2 => n17686, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_14_port, B2 => 
                           n14245, C1 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_14_port, C2 => 
                           n17687, ZN => n14590);
   U9066 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_27_14_port,
                           A2 => n17688, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_14_port, B2 => 
                           n17689, ZN => n14584);
   U9065 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_23_14_port,
                           A2 => n17690, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_14_port, B2 => 
                           n17691, ZN => n14585);
   U9064 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_21_14_port,
                           A2 => n17692, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_14_port, B2 => 
                           n17693, ZN => n14586);
   U9063 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_19_14_port,
                           A2 => n17694, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_14_port, B2 => 
                           n17695, ZN => n14587);
   U9062 : NAND4_X1 port map( A1 => n14584, A2 => n14585, A3 => n14586, A4 => 
                           n14587, ZN => n14573);
   U9061 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_17_14_port,
                           A2 => n17696, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_14_port, B2 => 
                           n17697, ZN => n14580);
   U9060 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_12_14_port,
                           A2 => n17698, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_14_port, B2 => 
                           n17358, ZN => n14581);
   U9059 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_8_14_port, 
                           A2 => n14223, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_14_port, B2 => 
                           n17152, ZN => n14582);
   U9058 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_9_14_port, 
                           A2 => n17352, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_14_port, B2 => 
                           n17699, ZN => n14583);
   U9057 : NAND4_X1 port map( A1 => n14580, A2 => n14581, A3 => n14582, A4 => 
                           n14583, ZN => n14574);
   U9056 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_11_14_port,
                           A2 => n14215, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_14_port, B2 => 
                           n14216, ZN => n14576);
   U9055 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_14_14_port,
                           A2 => n14213, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_14_port, B2 => 
                           n14214, ZN => n14577);
   U9054 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_2_14_port, 
                           A2 => n17355, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_14_port, B2 => 
                           n14212, ZN => n14578);
   U9053 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_6_14_port, 
                           A2 => n17356, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_14_port, B2 => 
                           n14210, ZN => n14579);
   U9052 : NAND4_X1 port map( A1 => n14576, A2 => n14577, A3 => n14578, A4 => 
                           n14579, ZN => n14575);
   U9051 : NOR4_X1 port map( A1 => n14572, A2 => n14573, A3 => n14574, A4 => 
                           n14575, ZN => n14571);
   U9050 : NOR2_X1 port map( A1 => n14571, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N148);
   U8729 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_31_31_port,
                           A2 => n14249, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_31_port, B2 => 
                           n14250, ZN => n14241);
   U8728 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_29_31_port,
                           A2 => n14247, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_31_port, B2 => 
                           n14248, ZN => n14242);
   U8727 : AOI222_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_4_31_port,
                           A2 => n14244, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_31_port, B2 => 
                           n14245, C1 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_31_port, C2 => 
                           n17687, ZN => n14243);
   U8726 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_27_31_port,
                           A2 => n14239, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_31_port, B2 => 
                           n14240, ZN => n14229);
   U8725 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_23_31_port,
                           A2 => n14237, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_31_port, B2 => 
                           n14238, ZN => n14230);
   U8724 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_21_31_port,
                           A2 => n14235, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_31_port, B2 => 
                           n14236, ZN => n14231);
   U8723 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_19_31_port,
                           A2 => n14233, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_31_port, B2 => 
                           n14234, ZN => n14232);
   U8722 : NAND4_X1 port map( A1 => n14229, A2 => n14230, A3 => n14231, A4 => 
                           n14232, ZN => n14202);
   U8721 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_17_31_port,
                           A2 => n14227, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_31_port, B2 => 
                           n14228, ZN => n14217);
   U8720 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_12_31_port,
                           A2 => n14225, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_31_port, B2 => 
                           n17358, ZN => n14218);
   U8719 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_8_31_port, 
                           A2 => n14223, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_31_port, B2 => 
                           n17152, ZN => n14219);
   U8718 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_9_31_port, 
                           A2 => n17352, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_31_port, B2 => 
                           n14222, ZN => n14220);
   U8717 : NAND4_X1 port map( A1 => n14217, A2 => n14218, A3 => n14219, A4 => 
                           n14220, ZN => n14203);
   U8716 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_11_31_port,
                           A2 => n17151, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_31_port, B2 => 
                           n14216, ZN => n14205);
   U8715 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_14_31_port,
                           A2 => n17700, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_31_port, B2 => 
                           n14214, ZN => n14206);
   U8714 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_2_31_port, 
                           A2 => n17355, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_31_port, B2 => 
                           n14212, ZN => n14207);
   U8713 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_6_31_port, 
                           A2 => n17356, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_31_port, B2 => 
                           n14210, ZN => n14208);
   U8712 : NAND4_X1 port map( A1 => n14205, A2 => n14206, A3 => n14207, A4 => 
                           n14208, ZN => n14204);
   U8711 : NOR4_X1 port map( A1 => n14201, A2 => n14202, A3 => n14203, A4 => 
                           n14204, ZN => n14200);
   U8710 : NOR2_X1 port map( A1 => n14200, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N165);
   U9149 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_31_10_port,
                           A2 => n17154, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_10_port, B2 => 
                           n17683, ZN => n14668);
   U9148 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_29_10_port,
                           A2 => n17684, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_10_port, B2 => 
                           n17685, ZN => n14669);
   U9147 : AOI222_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_4_10_port,
                           A2 => n17686, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_10_port, B2 => 
                           n17153, C1 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_10_port, C2 => 
                           n17687, ZN => n14670);
   U9146 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_27_10_port,
                           A2 => n17688, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_10_port, B2 => 
                           n17689, ZN => n14664);
   U9145 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_23_10_port,
                           A2 => n17690, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_10_port, B2 => 
                           n17691, ZN => n14665);
   U9144 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_21_10_port,
                           A2 => n17692, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_10_port, B2 => 
                           n17693, ZN => n14666);
   U9143 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_19_10_port,
                           A2 => n17694, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_10_port, B2 => 
                           n17695, ZN => n14667);
   U9142 : NAND4_X1 port map( A1 => n14664, A2 => n14665, A3 => n14666, A4 => 
                           n14667, ZN => n14653);
   U9141 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_17_10_port,
                           A2 => n17696, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_10_port, B2 => 
                           n17697, ZN => n14660);
   U9140 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_12_10_port,
                           A2 => n17698, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_10_port, B2 => 
                           n17358, ZN => n14661);
   U9139 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_8_10_port, 
                           A2 => n14223, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_10_port, B2 => 
                           n17152, ZN => n14662);
   U9138 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_9_10_port, 
                           A2 => n17352, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_10_port, B2 => 
                           n17699, ZN => n14663);
   U9137 : NAND4_X1 port map( A1 => n14660, A2 => n14661, A3 => n14662, A4 => 
                           n14663, ZN => n14654);
   U9136 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_11_10_port,
                           A2 => n17151, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_10_port, B2 => 
                           n14216, ZN => n14656);
   U9135 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_14_10_port,
                           A2 => n17700, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_10_port, B2 => 
                           n14214, ZN => n14657);
   U9134 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_2_10_port, 
                           A2 => n17355, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_10_port, B2 => 
                           n14212, ZN => n14658);
   U9133 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_6_10_port, 
                           A2 => n17356, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_10_port, B2 => 
                           n14210, ZN => n14659);
   U9132 : NAND4_X1 port map( A1 => n14656, A2 => n14657, A3 => n14658, A4 => 
                           n14659, ZN => n14655);
   U9131 : NOR4_X1 port map( A1 => n14652, A2 => n14653, A3 => n14654, A4 => 
                           n14655, ZN => n14651);
   U9130 : NOR2_X1 port map( A1 => n14651, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N144);
   U8829 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_31_26_port,
                           A2 => n17154, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_26_port, B2 => 
                           n17683, ZN => n14348);
   U8828 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_29_26_port,
                           A2 => n17684, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_26_port, B2 => 
                           n17685, ZN => n14349);
   U8827 : AOI222_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_4_26_port,
                           A2 => n17686, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_26_port, B2 => 
                           n17153, C1 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_26_port, C2 => 
                           n17687, ZN => n14350);
   U8826 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_27_26_port,
                           A2 => n17688, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_26_port, B2 => 
                           n17689, ZN => n14344);
   U8825 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_23_26_port,
                           A2 => n17690, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_26_port, B2 => 
                           n17691, ZN => n14345);
   U8824 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_21_26_port,
                           A2 => n17692, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_26_port, B2 => 
                           n17693, ZN => n14346);
   U8823 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_19_26_port,
                           A2 => n17694, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_26_port, B2 => 
                           n17695, ZN => n14347);
   U8822 : NAND4_X1 port map( A1 => n14344, A2 => n14345, A3 => n14346, A4 => 
                           n14347, ZN => n14333);
   U8821 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_17_26_port,
                           A2 => n17696, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_26_port, B2 => 
                           n17697, ZN => n14340);
   U8820 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_12_26_port,
                           A2 => n17698, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_26_port, B2 => 
                           n17357, ZN => n14341);
   U8819 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_8_26_port, 
                           A2 => n17417, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_26_port, B2 => 
                           n14224, ZN => n14342);
   U8818 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_9_26_port, 
                           A2 => n17351, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_26_port, B2 => 
                           n17699, ZN => n14343);
   U8817 : NAND4_X1 port map( A1 => n14340, A2 => n14341, A3 => n14342, A4 => 
                           n14343, ZN => n14334);
   U8816 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_11_26_port,
                           A2 => n17151, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_26_port, B2 => 
                           n17413, ZN => n14336);
   U8815 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_14_26_port,
                           A2 => n17700, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_26_port, B2 => 
                           n17414, ZN => n14337);
   U8814 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_2_26_port, 
                           A2 => n17353, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_26_port, B2 => 
                           n17415, ZN => n14338);
   U8813 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_6_26_port, 
                           A2 => n17354, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_26_port, B2 => 
                           n17416, ZN => n14339);
   U8812 : NAND4_X1 port map( A1 => n14336, A2 => n14337, A3 => n14338, A4 => 
                           n14339, ZN => n14335);
   U8811 : NOR4_X1 port map( A1 => n14332, A2 => n14333, A3 => n14334, A4 => 
                           n14335, ZN => n14331);
   U8810 : NOR2_X1 port map( A1 => n14331, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N160);
   U9329 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_31_1_port, 
                           A2 => n17154, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_1_port, B2 => 
                           n17683, ZN => n14848);
   U9328 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_29_1_port, 
                           A2 => n17684, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_1_port, B2 => 
                           n17685, ZN => n14849);
   U9327 : AOI222_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_4_1_port, 
                           A2 => n17686, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_1_port, B2 => 
                           n17153, C1 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_1_port, C2 => 
                           n17687, ZN => n14850);
   U9326 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_27_1_port, 
                           A2 => n17688, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_1_port, B2 => 
                           n17689, ZN => n14844);
   U9325 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_23_1_port, 
                           A2 => n17690, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_1_port, B2 => 
                           n17691, ZN => n14845);
   U9324 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_21_1_port, 
                           A2 => n17692, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_1_port, B2 => 
                           n17693, ZN => n14846);
   U9323 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_19_1_port, 
                           A2 => n17694, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_1_port, B2 => 
                           n17695, ZN => n14847);
   U9322 : NAND4_X1 port map( A1 => n14844, A2 => n14845, A3 => n14846, A4 => 
                           n14847, ZN => n14833);
   U9321 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_17_1_port, 
                           A2 => n17696, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_1_port, B2 => 
                           n17697, ZN => n14840);
   U9320 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_12_1_port, 
                           A2 => n17698, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_1_port, B2 => 
                           n17357, ZN => n14841);
   U9319 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_8_1_port, 
                           A2 => n17417, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_1_port, B2 => 
                           n14224, ZN => n14842);
   U9318 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_9_1_port, 
                           A2 => n17351, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_1_port, B2 => 
                           n17699, ZN => n14843);
   U9317 : NAND4_X1 port map( A1 => n14840, A2 => n14841, A3 => n14842, A4 => 
                           n14843, ZN => n14834);
   U9316 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_11_1_port, 
                           A2 => n17151, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_1_port, B2 => 
                           n17413, ZN => n14836);
   U9315 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_14_1_port, 
                           A2 => n17700, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_1_port, B2 => 
                           n17414, ZN => n14837);
   U9314 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_2_1_port, 
                           A2 => n17353, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_1_port, B2 => 
                           n17415, ZN => n14838);
   U9313 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_6_1_port, 
                           A2 => n17354, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_1_port, B2 => 
                           n17416, ZN => n14839);
   U9312 : NAND4_X1 port map( A1 => n14836, A2 => n14837, A3 => n14838, A4 => 
                           n14839, ZN => n14835);
   U9311 : NOR4_X1 port map( A1 => n14832, A2 => n14833, A3 => n14834, A4 => 
                           n14835, ZN => n14831);
   U9310 : NOR2_X1 port map( A1 => n14831, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N135);
   U8789 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_31_28_port,
                           A2 => n17154, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_28_port, B2 => 
                           n17683, ZN => n14308);
   U8788 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_29_28_port,
                           A2 => n17684, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_28_port, B2 => 
                           n17685, ZN => n14309);
   U8787 : AOI222_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_4_28_port,
                           A2 => n17686, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_28_port, B2 => 
                           n17153, C1 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_28_port, C2 => 
                           n17687, ZN => n14310);
   U8786 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_27_28_port,
                           A2 => n17688, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_28_port, B2 => 
                           n17689, ZN => n14304);
   U8785 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_23_28_port,
                           A2 => n17690, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_28_port, B2 => 
                           n17691, ZN => n14305);
   U8784 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_21_28_port,
                           A2 => n17692, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_28_port, B2 => 
                           n17693, ZN => n14306);
   U8783 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_19_28_port,
                           A2 => n17694, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_28_port, B2 => 
                           n17695, ZN => n14307);
   U8782 : NAND4_X1 port map( A1 => n14304, A2 => n14305, A3 => n14306, A4 => 
                           n14307, ZN => n14293);
   U8781 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_17_28_port,
                           A2 => n17696, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_28_port, B2 => 
                           n17697, ZN => n14300);
   U8780 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_12_28_port,
                           A2 => n17698, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_28_port, B2 => 
                           n17358, ZN => n14301);
   U8779 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_8_28_port, 
                           A2 => n17417, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_28_port, B2 => 
                           n14224, ZN => n14302);
   U8778 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_9_28_port, 
                           A2 => n17352, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_28_port, B2 => 
                           n17699, ZN => n14303);
   U8777 : NAND4_X1 port map( A1 => n14300, A2 => n14301, A3 => n14302, A4 => 
                           n14303, ZN => n14294);
   U8776 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_11_28_port,
                           A2 => n17151, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_28_port, B2 => 
                           n17413, ZN => n14296);
   U8775 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_14_28_port,
                           A2 => n17700, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_28_port, B2 => 
                           n17414, ZN => n14297);
   U8774 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_2_28_port, 
                           A2 => n17355, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_28_port, B2 => 
                           n17415, ZN => n14298);
   U8773 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_6_28_port, 
                           A2 => n17356, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_28_port, B2 => 
                           n17416, ZN => n14299);
   U8772 : NAND4_X1 port map( A1 => n14296, A2 => n14297, A3 => n14298, A4 => 
                           n14299, ZN => n14295);
   U8771 : NOR4_X1 port map( A1 => n14292, A2 => n14293, A3 => n14294, A4 => 
                           n14295, ZN => n14291);
   U8770 : NOR2_X1 port map( A1 => n14291, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N162);
   U9189 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_31_8_port, 
                           A2 => n17154, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_8_port, B2 => 
                           n17683, ZN => n14708);
   U9188 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_29_8_port, 
                           A2 => n17684, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_8_port, B2 => 
                           n17685, ZN => n14709);
   U9187 : AOI222_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_4_8_port, 
                           A2 => n17686, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_8_port, B2 => 
                           n17153, C1 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_8_port, C2 => 
                           n17687, ZN => n14710);
   U9186 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_27_8_port, 
                           A2 => n17688, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_8_port, B2 => 
                           n17689, ZN => n14704);
   U9185 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_23_8_port, 
                           A2 => n17690, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_8_port, B2 => 
                           n17691, ZN => n14705);
   U9184 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_21_8_port, 
                           A2 => n17692, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_8_port, B2 => 
                           n17693, ZN => n14706);
   U9183 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_19_8_port, 
                           A2 => n17694, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_8_port, B2 => 
                           n17695, ZN => n14707);
   U9182 : NAND4_X1 port map( A1 => n14704, A2 => n14705, A3 => n14706, A4 => 
                           n14707, ZN => n14693);
   U9181 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_17_8_port, 
                           A2 => n17696, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_8_port, B2 => 
                           n17697, ZN => n14700);
   U9180 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_12_8_port, 
                           A2 => n17698, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_8_port, B2 => 
                           n17358, ZN => n14701);
   U9179 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_8_8_port, 
                           A2 => n17417, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_8_port, B2 => 
                           n17152, ZN => n14702);
   U9178 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_9_8_port, 
                           A2 => n17352, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_8_port, B2 => 
                           n17699, ZN => n14703);
   U9177 : NAND4_X1 port map( A1 => n14700, A2 => n14701, A3 => n14702, A4 => 
                           n14703, ZN => n14694);
   U9176 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_11_8_port, 
                           A2 => n17151, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_8_port, B2 => 
                           n17413, ZN => n14696);
   U9175 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_14_8_port, 
                           A2 => n17700, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_8_port, B2 => 
                           n17414, ZN => n14697);
   U9174 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_2_8_port, 
                           A2 => n17355, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_8_port, B2 => 
                           n17415, ZN => n14698);
   U9173 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_6_8_port, 
                           A2 => n17356, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_8_port, B2 => 
                           n17416, ZN => n14699);
   U9172 : NAND4_X1 port map( A1 => n14696, A2 => n14697, A3 => n14698, A4 => 
                           n14699, ZN => n14695);
   U9171 : NOR4_X1 port map( A1 => n14692, A2 => n14693, A3 => n14694, A4 => 
                           n14695, ZN => n14691);
   U9170 : NOR2_X1 port map( A1 => n14691, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N142);
   U8869 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_31_24_port,
                           A2 => n17154, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_24_port, B2 => 
                           n17683, ZN => n14388);
   U8868 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_29_24_port,
                           A2 => n17684, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_24_port, B2 => 
                           n17685, ZN => n14389);
   U8867 : AOI222_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_4_24_port,
                           A2 => n17686, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_24_port, B2 => 
                           n17153, C1 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_24_port, C2 => 
                           n17687, ZN => n14390);
   U8866 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_27_24_port,
                           A2 => n17688, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_24_port, B2 => 
                           n17689, ZN => n14384);
   U8865 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_23_24_port,
                           A2 => n17690, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_24_port, B2 => 
                           n17691, ZN => n14385);
   U8864 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_21_24_port,
                           A2 => n17692, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_24_port, B2 => 
                           n17693, ZN => n14386);
   U8863 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_19_24_port,
                           A2 => n17694, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_24_port, B2 => 
                           n17695, ZN => n14387);
   U8862 : NAND4_X1 port map( A1 => n14384, A2 => n14385, A3 => n14386, A4 => 
                           n14387, ZN => n14373);
   U8861 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_17_24_port,
                           A2 => n17696, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_24_port, B2 => 
                           n17697, ZN => n14380);
   U8860 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_12_24_port,
                           A2 => n17698, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_24_port, B2 => 
                           n17357, ZN => n14381);
   U8859 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_8_24_port, 
                           A2 => n17417, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_24_port, B2 => 
                           n14224, ZN => n14382);
   U8858 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_9_24_port, 
                           A2 => n17351, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_24_port, B2 => 
                           n17699, ZN => n14383);
   U8857 : NAND4_X1 port map( A1 => n14380, A2 => n14381, A3 => n14382, A4 => 
                           n14383, ZN => n14374);
   U8856 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_11_24_port,
                           A2 => n17151, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_24_port, B2 => 
                           n17413, ZN => n14376);
   U8855 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_14_24_port,
                           A2 => n17700, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_24_port, B2 => 
                           n17414, ZN => n14377);
   U8854 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_2_24_port, 
                           A2 => n17353, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_24_port, B2 => 
                           n17415, ZN => n14378);
   U8853 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_6_24_port, 
                           A2 => n17354, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_24_port, B2 => 
                           n17416, ZN => n14379);
   U8852 : NAND4_X1 port map( A1 => n14376, A2 => n14377, A3 => n14378, A4 => 
                           n14379, ZN => n14375);
   U8851 : NOR4_X1 port map( A1 => n14372, A2 => n14373, A3 => n14374, A4 => 
                           n14375, ZN => n14371);
   U8850 : NOR2_X1 port map( A1 => n14371, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N158);
   U9309 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_31_2_port, 
                           A2 => n17154, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_2_port, B2 => 
                           n17683, ZN => n14828);
   U9308 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_29_2_port, 
                           A2 => n17684, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_2_port, B2 => 
                           n17685, ZN => n14829);
   U9307 : AOI222_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_4_2_port, 
                           A2 => n14244, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_2_port, B2 => 
                           n17153, C1 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_2_port, C2 => 
                           n14246, ZN => n14830);
   U9306 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_27_2_port, 
                           A2 => n17688, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_2_port, B2 => 
                           n14240, ZN => n14824);
   U9305 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_23_2_port, 
                           A2 => n17690, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_2_port, B2 => 
                           n17691, ZN => n14825);
   U9304 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_21_2_port, 
                           A2 => n17692, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_2_port, B2 => 
                           n14236, ZN => n14826);
   U9303 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_19_2_port, 
                           A2 => n17694, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_2_port, B2 => 
                           n17695, ZN => n14827);
   U9302 : NAND4_X1 port map( A1 => n14824, A2 => n14825, A3 => n14826, A4 => 
                           n14827, ZN => n14813);
   U9301 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_17_2_port, 
                           A2 => n17696, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_2_port, B2 => 
                           n14228, ZN => n14820);
   U9300 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_12_2_port, 
                           A2 => n17698, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_2_port, B2 => 
                           n17357, ZN => n14821);
   U9299 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_8_2_port, 
                           A2 => n17417, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_2_port, B2 => 
                           n17152, ZN => n14822);
   U9298 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_9_2_port, 
                           A2 => n17351, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_2_port, B2 => 
                           n17699, ZN => n14823);
   U9297 : NAND4_X1 port map( A1 => n14820, A2 => n14821, A3 => n14822, A4 => 
                           n14823, ZN => n14814);
   U9296 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_11_2_port, 
                           A2 => n17151, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_2_port, B2 => 
                           n17413, ZN => n14816);
   U9295 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_14_2_port, 
                           A2 => n17700, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_2_port, B2 => 
                           n17414, ZN => n14817);
   U9294 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_2_2_port, 
                           A2 => n17353, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_2_port, B2 => 
                           n17415, ZN => n14818);
   U9293 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_6_2_port, 
                           A2 => n17354, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_2_port, B2 => 
                           n17416, ZN => n14819);
   U9292 : NAND4_X1 port map( A1 => n14816, A2 => n14817, A3 => n14818, A4 => 
                           n14819, ZN => n14815);
   U9291 : NOR4_X1 port map( A1 => n14812, A2 => n14813, A3 => n14814, A4 => 
                           n14815, ZN => n14811);
   U9290 : AOI21_X1 port map( B1 => n14025, B2 => n14811, A => n14168, ZN => 
                           pipeline_IDEX_Stage_N136);
   U8655 : NOR2_X1 port map( A1 => n17313, A2 => n14059, ZN => n14084);
   U8653 : NAND2_X1 port map( A1 => pipeline_inst_IFID_DEC_29_port, A2 => 
                           n14190, ZN => n13998);
   U8651 : NOR2_X1 port map( A1 => n17347, A2 => n14058, ZN => n13999);
   U8650 : NAND2_X1 port map( A1 => pipeline_inst_IFID_DEC_30_port, A2 => 
                           pipeline_inst_IFID_DEC_26_port, ZN => n14189);
   U8649 : NOR4_X1 port map( A1 => pipeline_inst_IFID_DEC_27_port, A2 => n17382
                           , A3 => n17348, A4 => n14189, ZN => n14040);
   U8648 : NOR2_X1 port map( A1 => n13999, A2 => n14040, ZN => n14042);
   U8647 : NAND2_X1 port map( A1 => n17313, A2 => n14001, ZN => n14011);
   U8645 : NAND2_X1 port map( A1 => pipeline_inst_IFID_DEC_30_port, A2 => 
                           n14185, ZN => n13997);
   U8644 : NAND2_X1 port map( A1 => n14042, A2 => n13997, ZN => n14016);
   U8643 : NOR4_X1 port map( A1 => n17313, A2 => n17347, A3 => n17382, A4 => 
                           pipeline_inst_IFID_DEC_28_port, ZN => n14022);
   U8642 : NOR2_X1 port map( A1 => n14016, A2 => n14022, ZN => n14188);
   U8641 : NAND2_X1 port map( A1 => n14029, A2 => n14188, ZN => n14009);
   U8640 : NAND2_X1 port map( A1 => n14049, A2 => 
                           pipeline_inst_IFID_DEC_29_port, ZN => n14187);
   U8639 : AOI21_X1 port map( B1 => pipeline_inst_IFID_DEC_27_port, B2 => 
                           n14176, A => n14187, ZN => n14183);
   U8638 : NAND2_X1 port map( A1 => pipeline_inst_IFID_DEC_30_port, A2 => 
                           n17409, ZN => n14047);
   U8637 : NOR2_X1 port map( A1 => n14186, A2 => n14047, ZN => n14061);
   U8636 : AOI21_X1 port map( B1 => n14185, B2 => n17347, A => n14061, ZN => 
                           n14028);
   U8635 : NAND4_X1 port map( A1 => n14049, A2 => n17382, A3 => 
                           pipeline_inst_IFID_DEC_27_port, A4 => 
                           pipeline_inst_IFID_DEC_30_port, ZN => n14019);
   U8634 : NAND2_X1 port map( A1 => n14028, A2 => n14019, ZN => n14184);
   U8632 : NAND2_X1 port map( A1 => pipeline_stageD_offset_to_jump_temp_5_port,
                           A2 => n17404, ZN => n14181);
   U8631 : NOR3_X1 port map( A1 => pipeline_stageD_offset_to_jump_temp_4_port, 
                           A2 => pipeline_stageD_offset_to_jump_temp_3_port, A3
                           => n17404, ZN => n14067);
   U8628 : NAND2_X1 port map( A1 => n14179, A2 => n14051, ZN => n14024);
   U8627 : OAI211_X1 port map( C1 => pipeline_stageD_offset_to_jump_temp_4_port
                           , C2 => n14181, A => n14066, B => n14024, ZN => 
                           n14172);
   U8625 : NOR2_X1 port map( A1 => n17406, A2 => n17076, ZN => n14031);
   U8624 : OAI221_X1 port map( B1 => n14032, B2 => n14031, C1 => n14032, C2 => 
                           n17350, A => n14067, ZN => n14178);
   U8621 : NOR2_X1 port map( A1 => pipeline_stageD_offset_to_jump_temp_4_port, 
                           A2 => n14180, ZN => n14065);
   U8619 : NOR2_X1 port map( A1 => n17076, A2 => n14180, ZN => n14045);
   U8618 : AOI21_X1 port map( B1 => n14031, B2 => n14179, A => n14045, ZN => 
                           n14023);
   U8617 : NAND2_X1 port map( A1 => n14051, A2 => n14067, ZN => n14064);
   U8616 : NAND4_X1 port map( A1 => n14178, A2 => n14006, A3 => n14023, A4 => 
                           n14064, ZN => n14173);
   U8613 : OAI21_X1 port map( B1 => n14172, B2 => n14173, A => n14005, ZN => 
                           n14170);
   U8612 : OAI221_X1 port map( B1 => n14168, B2 => n13980, C1 => n14168, C2 => 
                           n14170, A => n17682, ZN => pipeline_IDEX_Stage_N90);
   U9438 : OAI22_X1 port map( A1 => n14931, A2 => n17075, B1 => n17109, B2 => 
                           n17468, ZN => pipeline_IDEX_Stage_N109);
   U9430 : OAI22_X1 port map( A1 => n14923, A2 => n17075, B1 => n17682, B2 => 
                           n17441, ZN => pipeline_IDEX_Stage_N113);
   U9412 : OAI22_X1 port map( A1 => n14905, A2 => n17075, B1 => n17682, B2 => 
                           n17463, ZN => pipeline_IDEX_Stage_N122);
   U9446 : OAI22_X1 port map( A1 => n14939, A2 => n17075, B1 => n17109, B2 => 
                           n17439, ZN => pipeline_IDEX_Stage_N105);
   U9428 : OAI22_X1 port map( A1 => n14921, A2 => n17075, B1 => n17109, B2 => 
                           n17459, ZN => pipeline_IDEX_Stage_N114);
   U9436 : OAI22_X1 port map( A1 => n14929, A2 => n17075, B1 => n17109, B2 => 
                           n17457, ZN => pipeline_IDEX_Stage_N110);
   U9410 : OAI22_X1 port map( A1 => n14903, A2 => n17075, B1 => n17109, B2 => 
                           n17448, ZN => pipeline_IDEX_Stage_N123);
   U9418 : OAI22_X1 port map( A1 => n14911, A2 => n17075, B1 => n17109, B2 => 
                           n17443, ZN => pipeline_IDEX_Stage_N119);
   U9444 : OAI22_X1 port map( A1 => n14937, A2 => n17075, B1 => n17109, B2 => 
                           n17455, ZN => pipeline_IDEX_Stage_N106);
   U9400 : OAI22_X1 port map( A1 => n14893, A2 => n17075, B1 => n17682, B2 => 
                           n17466, ZN => pipeline_IDEX_Stage_N128);
   U9440 : OAI22_X1 port map( A1 => n14933, A2 => n17075, B1 => n17682, B2 => 
                           n17456, ZN => pipeline_IDEX_Stage_N108);
   U9398 : OAI22_X1 port map( A1 => n14891, A2 => n17075, B1 => n17682, B2 => 
                           n17469, ZN => pipeline_IDEX_Stage_N129);
   U9450 : OAI22_X1 port map( A1 => n14943, A2 => n17075, B1 => n17109, B2 => 
                           n17446, ZN => pipeline_IDEX_Stage_N103);
   U9406 : OAI22_X1 port map( A1 => n14899, A2 => n17075, B1 => n17682, B2 => 
                           n17435, ZN => pipeline_IDEX_Stage_N125);
   U9404 : OAI22_X1 port map( A1 => n14897, A2 => n17075, B1 => n17682, B2 => 
                           n17465, ZN => pipeline_IDEX_Stage_N126);
   U9448 : OAI22_X1 port map( A1 => n14941, A2 => n17075, B1 => n17682, B2 => 
                           n17470, ZN => pipeline_IDEX_Stage_N104);
   U9396 : OAI22_X1 port map( A1 => n14889, A2 => n17075, B1 => n17109, B2 => 
                           n17467, ZN => pipeline_IDEX_Stage_N130);
   U9434 : OAI22_X1 port map( A1 => n14927, A2 => n17075, B1 => n17109, B2 => 
                           n17436, ZN => pipeline_IDEX_Stage_N111);
   U9426 : OAI22_X1 port map( A1 => n14919, A2 => n17075, B1 => n17109, B2 => 
                           n17442, ZN => pipeline_IDEX_Stage_N115);
   U9392 : OAI22_X1 port map( A1 => n14885, A2 => n17075, B1 => n17109, B2 => 
                           n17471, ZN => pipeline_IDEX_Stage_N132);
   U9432 : OAI22_X1 port map( A1 => n14925, A2 => n17075, B1 => n17109, B2 => 
                           n17458, ZN => pipeline_IDEX_Stage_N112);
   U9416 : OAI22_X1 port map( A1 => n14909, A2 => n17075, B1 => n17109, B2 => 
                           n17462, ZN => pipeline_IDEX_Stage_N120);
   U9408 : OAI22_X1 port map( A1 => n14901, A2 => n17075, B1 => n17109, B2 => 
                           n17464, ZN => pipeline_IDEX_Stage_N124);
   U8949 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_31_20_port,
                           A2 => n17154, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_20_port, B2 => 
                           n17683, ZN => n14468);
   U8948 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_29_20_port,
                           A2 => n17684, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_20_port, B2 => 
                           n17685, ZN => n14469);
   U8947 : AOI222_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_4_20_port,
                           A2 => n14244, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_20_port, B2 => 
                           n17153, C1 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_20_port, C2 => 
                           n14246, ZN => n14470);
   U8946 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_27_20_port,
                           A2 => n17688, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_20_port, B2 => 
                           n14240, ZN => n14464);
   U8945 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_23_20_port,
                           A2 => n17690, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_20_port, B2 => 
                           n17691, ZN => n14465);
   U8944 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_21_20_port,
                           A2 => n17692, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_20_port, B2 => 
                           n14236, ZN => n14466);
   U8943 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_19_20_port,
                           A2 => n17694, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_20_port, B2 => 
                           n17695, ZN => n14467);
   U8942 : NAND4_X1 port map( A1 => n14464, A2 => n14465, A3 => n14466, A4 => 
                           n14467, ZN => n14453);
   U8941 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_17_20_port,
                           A2 => n17696, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_20_port, B2 => 
                           n14228, ZN => n14460);
   U8940 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_12_20_port,
                           A2 => n17698, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_20_port, B2 => 
                           n14226, ZN => n14461);
   U8939 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_8_20_port, 
                           A2 => n14223, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_20_port, B2 => 
                           n17152, ZN => n14462);
   U8938 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_9_20_port, 
                           A2 => n14221, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_20_port, B2 => 
                           n17699, ZN => n14463);
   U8937 : NAND4_X1 port map( A1 => n14460, A2 => n14461, A3 => n14462, A4 => 
                           n14463, ZN => n14454);
   U8936 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_11_20_port,
                           A2 => n17151, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_20_port, B2 => 
                           n14216, ZN => n14456);
   U8935 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_14_20_port,
                           A2 => n17700, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_20_port, B2 => 
                           n14214, ZN => n14457);
   U8934 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_2_20_port, 
                           A2 => n17367, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_20_port, B2 => 
                           n14212, ZN => n14458);
   U8933 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_6_20_port, 
                           A2 => n17368, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_20_port, B2 => 
                           n14210, ZN => n14459);
   U8932 : NAND4_X1 port map( A1 => n14456, A2 => n14457, A3 => n14458, A4 => 
                           n14459, ZN => n14455);
   U8931 : NOR4_X1 port map( A1 => n14452, A2 => n14453, A3 => n14454, A4 => 
                           n14455, ZN => n14451);
   U8930 : NOR2_X1 port map( A1 => n14451, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N154);
   U8929 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_31_21_port,
                           A2 => n17154, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_21_port, B2 => 
                           n14250, ZN => n14448);
   U8928 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_29_21_port,
                           A2 => n17684, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_21_port, B2 => 
                           n14248, ZN => n14449);
   U8927 : AOI222_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_4_21_port,
                           A2 => n17686, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_21_port, B2 => 
                           n17153, C1 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_21_port, C2 => 
                           n17687, ZN => n14450);
   U8926 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_27_21_port,
                           A2 => n17688, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_21_port, B2 => 
                           n17689, ZN => n14444);
   U8925 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_23_21_port,
                           A2 => n17690, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_21_port, B2 => 
                           n14238, ZN => n14445);
   U8924 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_21_21_port,
                           A2 => n14235, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_21_port, B2 => 
                           n17693, ZN => n14446);
   U8923 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_19_21_port,
                           A2 => n14233, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_21_port, B2 => 
                           n17695, ZN => n14447);
   U8922 : NAND4_X1 port map( A1 => n14444, A2 => n14445, A3 => n14446, A4 => 
                           n14447, ZN => n14433);
   U8921 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_17_21_port,
                           A2 => n17696, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_21_port, B2 => 
                           n17697, ZN => n14440);
   U8920 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_12_21_port,
                           A2 => n14225, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_21_port, B2 => 
                           n14226, ZN => n14441);
   U8919 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_8_21_port, 
                           A2 => n14223, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_21_port, B2 => 
                           n17152, ZN => n14442);
   U8918 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_9_21_port, 
                           A2 => n14221, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_21_port, B2 => 
                           n17699, ZN => n14443);
   U8917 : NAND4_X1 port map( A1 => n14440, A2 => n14441, A3 => n14442, A4 => 
                           n14443, ZN => n14434);
   U8916 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_11_21_port,
                           A2 => n17151, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_21_port, B2 => 
                           n14216, ZN => n14436);
   U8915 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_14_21_port,
                           A2 => n14213, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_21_port, B2 => 
                           n14214, ZN => n14437);
   U8914 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_2_21_port, 
                           A2 => n17367, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_21_port, B2 => 
                           n14212, ZN => n14438);
   U8913 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_6_21_port, 
                           A2 => n17368, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_21_port, B2 => 
                           n14210, ZN => n14439);
   U8912 : NAND4_X1 port map( A1 => n14436, A2 => n14437, A3 => n14438, A4 => 
                           n14439, ZN => n14435);
   U8911 : NOR4_X1 port map( A1 => n14432, A2 => n14433, A3 => n14434, A4 => 
                           n14435, ZN => n14431);
   U8910 : NOR2_X1 port map( A1 => n14431, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N155);
   U9029 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_31_16_port,
                           A2 => n17154, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_16_port, B2 => 
                           n14250, ZN => n14548);
   U9028 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_29_16_port,
                           A2 => n17684, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_16_port, B2 => 
                           n14248, ZN => n14549);
   U9027 : AOI222_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_4_16_port,
                           A2 => n14244, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_16_port, B2 => 
                           n17153, C1 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_16_port, C2 => 
                           n17687, ZN => n14550);
   U9026 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_27_16_port,
                           A2 => n17688, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_16_port, B2 => 
                           n14240, ZN => n14544);
   U9025 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_23_16_port,
                           A2 => n17690, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_16_port, B2 => 
                           n14238, ZN => n14545);
   U9024 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_21_16_port,
                           A2 => n17692, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_16_port, B2 => 
                           n14236, ZN => n14546);
   U9023 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_19_16_port,
                           A2 => n17694, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_16_port, B2 => 
                           n14234, ZN => n14547);
   U9022 : NAND4_X1 port map( A1 => n14544, A2 => n14545, A3 => n14546, A4 => 
                           n14547, ZN => n14533);
   U9021 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_17_16_port,
                           A2 => n17696, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_16_port, B2 => 
                           n14228, ZN => n14540);
   U9020 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_12_16_port,
                           A2 => n14225, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_16_port, B2 => 
                           n14226, ZN => n14541);
   U9019 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_8_16_port, 
                           A2 => n14223, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_16_port, B2 => 
                           n17152, ZN => n14542);
   U9018 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_9_16_port, 
                           A2 => n14221, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_16_port, B2 => 
                           n14222, ZN => n14543);
   U9017 : NAND4_X1 port map( A1 => n14540, A2 => n14541, A3 => n14542, A4 => 
                           n14543, ZN => n14534);
   U9016 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_11_16_port,
                           A2 => n17151, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_16_port, B2 => 
                           n14216, ZN => n14536);
   U9015 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_14_16_port,
                           A2 => n14213, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_16_port, B2 => 
                           n14214, ZN => n14537);
   U9014 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_2_16_port, 
                           A2 => n17367, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_16_port, B2 => 
                           n14212, ZN => n14538);
   U9013 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_6_16_port, 
                           A2 => n17368, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_16_port, B2 => 
                           n14210, ZN => n14539);
   U9012 : NAND4_X1 port map( A1 => n14536, A2 => n14537, A3 => n14538, A4 => 
                           n14539, ZN => n14535);
   U9011 : NOR4_X1 port map( A1 => n14532, A2 => n14533, A3 => n14534, A4 => 
                           n14535, ZN => n14531);
   U9010 : NOR2_X1 port map( A1 => n14531, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N150);
   U9109 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_31_12_port,
                           A2 => n17154, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_12_port, B2 => 
                           n14250, ZN => n14628);
   U9108 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_29_12_port,
                           A2 => n17684, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_12_port, B2 => 
                           n14248, ZN => n14629);
   U9107 : AOI222_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_4_12_port,
                           A2 => n17686, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_12_port, B2 => 
                           n17153, C1 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_12_port, C2 => 
                           n14246, ZN => n14630);
   U9106 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_27_12_port,
                           A2 => n14239, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_12_port, B2 => 
                           n17689, ZN => n14624);
   U9105 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_23_12_port,
                           A2 => n17690, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_12_port, B2 => 
                           n14238, ZN => n14625);
   U9104 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_21_12_port,
                           A2 => n17692, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_12_port, B2 => 
                           n17693, ZN => n14626);
   U9103 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_19_12_port,
                           A2 => n17694, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_12_port, B2 => 
                           n14234, ZN => n14627);
   U9102 : NAND4_X1 port map( A1 => n14624, A2 => n14625, A3 => n14626, A4 => 
                           n14627, ZN => n14613);
   U9101 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_17_12_port,
                           A2 => n14227, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_12_port, B2 => 
                           n17697, ZN => n14620);
   U9100 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_12_12_port,
                           A2 => n17698, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_12_port, B2 => 
                           n14226, ZN => n14621);
   U9099 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_8_12_port, 
                           A2 => n14223, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_12_port, B2 => 
                           n17152, ZN => n14622);
   U9098 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_9_12_port, 
                           A2 => n14221, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_12_port, B2 => 
                           n14222, ZN => n14623);
   U9097 : NAND4_X1 port map( A1 => n14620, A2 => n14621, A3 => n14622, A4 => 
                           n14623, ZN => n14614);
   U9096 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_11_12_port,
                           A2 => n17151, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_12_port, B2 => 
                           n14216, ZN => n14616);
   U9095 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_14_12_port,
                           A2 => n14213, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_12_port, B2 => 
                           n14214, ZN => n14617);
   U9094 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_2_12_port, 
                           A2 => n17367, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_12_port, B2 => 
                           n14212, ZN => n14618);
   U9093 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_6_12_port, 
                           A2 => n17368, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_12_port, B2 => 
                           n14210, ZN => n14619);
   U9092 : NAND4_X1 port map( A1 => n14616, A2 => n14617, A3 => n14618, A4 => 
                           n14619, ZN => n14615);
   U9091 : NOR4_X1 port map( A1 => n14612, A2 => n14613, A3 => n14614, A4 => 
                           n14615, ZN => n14611);
   U9090 : NOR2_X1 port map( A1 => n14611, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N146);
   U9209 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_31_7_port, 
                           A2 => n17154, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_7_port, B2 => 
                           n17683, ZN => n14728);
   U9208 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_29_7_port, 
                           A2 => n17684, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_7_port, B2 => 
                           n17685, ZN => n14729);
   U9207 : AOI222_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_4_7_port, 
                           A2 => n17686, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_7_port, B2 => 
                           n17153, C1 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_7_port, C2 => 
                           n17687, ZN => n14730);
   U9206 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_27_7_port, 
                           A2 => n17688, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_7_port, B2 => 
                           n17689, ZN => n14724);
   U9205 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_23_7_port, 
                           A2 => n17690, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_7_port, B2 => 
                           n17691, ZN => n14725);
   U9204 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_21_7_port, 
                           A2 => n14235, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_7_port, B2 => 
                           n17693, ZN => n14726);
   U9203 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_19_7_port, 
                           A2 => n17694, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_7_port, B2 => 
                           n14234, ZN => n14727);
   U9202 : NAND4_X1 port map( A1 => n14724, A2 => n14725, A3 => n14726, A4 => 
                           n14727, ZN => n14713);
   U9201 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_17_7_port, 
                           A2 => n17696, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_7_port, B2 => 
                           n17697, ZN => n14720);
   U9200 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_12_7_port, 
                           A2 => n14225, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_7_port, B2 => 
                           n17358, ZN => n14721);
   U9199 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_8_7_port, 
                           A2 => n17417, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_7_port, B2 => 
                           n17152, ZN => n14722);
   U9198 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_9_7_port, 
                           A2 => n17352, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_7_port, B2 => 
                           n14222, ZN => n14723);
   U9197 : NAND4_X1 port map( A1 => n14720, A2 => n14721, A3 => n14722, A4 => 
                           n14723, ZN => n14714);
   U9196 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_11_7_port, 
                           A2 => n17151, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_7_port, B2 => 
                           n17413, ZN => n14716);
   U9195 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_14_7_port, 
                           A2 => n17700, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_7_port, B2 => 
                           n17414, ZN => n14717);
   U9194 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_2_7_port, 
                           A2 => n17355, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_7_port, B2 => 
                           n17415, ZN => n14718);
   U9193 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_6_7_port, 
                           A2 => n17356, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_7_port, B2 => 
                           n17416, ZN => n14719);
   U9192 : NAND4_X1 port map( A1 => n14716, A2 => n14717, A3 => n14718, A4 => 
                           n14719, ZN => n14715);
   U9191 : NOR4_X1 port map( A1 => n14712, A2 => n14713, A3 => n14714, A4 => 
                           n14715, ZN => n14711);
   U9190 : NOR2_X1 port map( A1 => n14711, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N141);
   U9129 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_31_11_port,
                           A2 => n17154, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_11_port, B2 => 
                           n17683, ZN => n14648);
   U9128 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_29_11_port,
                           A2 => n14247, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_11_port, B2 => 
                           n17685, ZN => n14649);
   U9127 : AOI222_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_4_11_port,
                           A2 => n17686, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_11_port, B2 => 
                           n17153, C1 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_11_port, C2 => 
                           n17687, ZN => n14650);
   U9126 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_27_11_port,
                           A2 => n17688, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_11_port, B2 => 
                           n17689, ZN => n14644);
   U9125 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_23_11_port,
                           A2 => n14237, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_11_port, B2 => 
                           n17691, ZN => n14645);
   U9124 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_21_11_port,
                           A2 => n17692, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_11_port, B2 => 
                           n17693, ZN => n14646);
   U9123 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_19_11_port,
                           A2 => n14233, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_11_port, B2 => 
                           n17695, ZN => n14647);
   U9122 : NAND4_X1 port map( A1 => n14644, A2 => n14645, A3 => n14646, A4 => 
                           n14647, ZN => n14633);
   U9121 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_17_11_port,
                           A2 => n17696, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_11_port, B2 => 
                           n17697, ZN => n14640);
   U9120 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_12_11_port,
                           A2 => n17698, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_11_port, B2 => 
                           n17358, ZN => n14641);
   U9119 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_8_11_port, 
                           A2 => n14223, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_11_port, B2 => 
                           n17152, ZN => n14642);
   U9118 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_9_11_port, 
                           A2 => n17352, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_11_port, B2 => 
                           n17699, ZN => n14643);
   U9117 : NAND4_X1 port map( A1 => n14640, A2 => n14641, A3 => n14642, A4 => 
                           n14643, ZN => n14634);
   U9116 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_11_11_port,
                           A2 => n17151, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_11_port, B2 => 
                           n14216, ZN => n14636);
   U9115 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_14_11_port,
                           A2 => n17700, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_11_port, B2 => 
                           n14214, ZN => n14637);
   U9114 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_2_11_port, 
                           A2 => n17355, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_11_port, B2 => 
                           n14212, ZN => n14638);
   U9113 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_6_11_port, 
                           A2 => n17356, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_11_port, B2 => 
                           n14210, ZN => n14639);
   U9112 : NAND4_X1 port map( A1 => n14636, A2 => n14637, A3 => n14638, A4 => 
                           n14639, ZN => n14635);
   U9111 : NOR4_X1 port map( A1 => n14632, A2 => n14633, A3 => n14634, A4 => 
                           n14635, ZN => n14631);
   U9110 : NOR2_X1 port map( A1 => n14631, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N145);
   U8769 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_31_29_port,
                           A2 => n17154, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_29_port, B2 => 
                           n17683, ZN => n14288);
   U8768 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_29_29_port,
                           A2 => n17684, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_29_port, B2 => 
                           n17685, ZN => n14289);
   U8767 : AOI222_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_4_29_port,
                           A2 => n17686, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_29_port, B2 => 
                           n17153, C1 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_29_port, C2 => 
                           n17687, ZN => n14290);
   U8766 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_27_29_port,
                           A2 => n17688, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_29_port, B2 => 
                           n17689, ZN => n14284);
   U8765 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_23_29_port,
                           A2 => n14237, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_29_port, B2 => 
                           n17691, ZN => n14285);
   U8764 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_21_29_port,
                           A2 => n17692, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_29_port, B2 => 
                           n17693, ZN => n14286);
   U8763 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_19_29_port,
                           A2 => n17694, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_29_port, B2 => 
                           n17695, ZN => n14287);
   U8762 : NAND4_X1 port map( A1 => n14284, A2 => n14285, A3 => n14286, A4 => 
                           n14287, ZN => n14273);
   U8761 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_17_29_port,
                           A2 => n17696, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_29_port, B2 => 
                           n17697, ZN => n14280);
   U8760 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_12_29_port,
                           A2 => n17698, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_29_port, B2 => 
                           n17358, ZN => n14281);
   U8759 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_8_29_port, 
                           A2 => n17417, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_29_port, B2 => 
                           n17152, ZN => n14282);
   U8758 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_9_29_port, 
                           A2 => n17352, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_29_port, B2 => 
                           n17699, ZN => n14283);
   U8757 : NAND4_X1 port map( A1 => n14280, A2 => n14281, A3 => n14282, A4 => 
                           n14283, ZN => n14274);
   U8756 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_11_29_port,
                           A2 => n17151, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_29_port, B2 => 
                           n17413, ZN => n14276);
   U8755 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_14_29_port,
                           A2 => n17700, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_29_port, B2 => 
                           n17414, ZN => n14277);
   U8754 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_2_29_port, 
                           A2 => n17355, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_29_port, B2 => 
                           n17415, ZN => n14278);
   U8753 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_6_29_port, 
                           A2 => n17356, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_29_port, B2 => 
                           n17416, ZN => n14279);
   U8752 : NAND4_X1 port map( A1 => n14276, A2 => n14277, A3 => n14278, A4 => 
                           n14279, ZN => n14275);
   U8751 : NOR4_X1 port map( A1 => n14272, A2 => n14273, A3 => n14274, A4 => 
                           n14275, ZN => n14271);
   U8750 : NOR2_X1 port map( A1 => n14271, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N163);
   U8749 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_31_30_port,
                           A2 => n17154, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_30_port, B2 => 
                           n17683, ZN => n14268);
   U8748 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_29_30_port,
                           A2 => n14247, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_30_port, B2 => 
                           n17685, ZN => n14269);
   U8747 : AOI222_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_4_30_port,
                           A2 => n17686, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_30_port, B2 => 
                           n17153, C1 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_30_port, C2 => 
                           n17687, ZN => n14270);
   U8746 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_27_30_port,
                           A2 => n17688, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_30_port, B2 => 
                           n17689, ZN => n14264);
   U8745 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_23_30_port,
                           A2 => n17690, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_30_port, B2 => 
                           n17691, ZN => n14265);
   U8744 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_21_30_port,
                           A2 => n17692, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_30_port, B2 => 
                           n17693, ZN => n14266);
   U8743 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_19_30_port,
                           A2 => n17694, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_30_port, B2 => 
                           n17695, ZN => n14267);
   U8742 : NAND4_X1 port map( A1 => n14264, A2 => n14265, A3 => n14266, A4 => 
                           n14267, ZN => n14253);
   U8741 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_17_30_port,
                           A2 => n17696, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_30_port, B2 => 
                           n17697, ZN => n14260);
   U8740 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_12_30_port,
                           A2 => n17698, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_30_port, B2 => 
                           n17358, ZN => n14261);
   U8739 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_8_30_port, 
                           A2 => n17417, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_30_port, B2 => 
                           n17152, ZN => n14262);
   U8738 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_9_30_port, 
                           A2 => n17352, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_30_port, B2 => 
                           n17699, ZN => n14263);
   U8737 : NAND4_X1 port map( A1 => n14260, A2 => n14261, A3 => n14262, A4 => 
                           n14263, ZN => n14254);
   U8736 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_11_30_port,
                           A2 => n17151, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_30_port, B2 => 
                           n17413, ZN => n14256);
   U8735 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_14_30_port,
                           A2 => n17700, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_30_port, B2 => 
                           n17414, ZN => n14257);
   U8734 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_2_30_port, 
                           A2 => n17355, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_30_port, B2 => 
                           n17415, ZN => n14258);
   U8733 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_6_30_port, 
                           A2 => n17356, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_30_port, B2 => 
                           n17416, ZN => n14259);
   U8732 : NAND4_X1 port map( A1 => n14256, A2 => n14257, A3 => n14258, A4 => 
                           n14259, ZN => n14255);
   U8731 : NOR4_X1 port map( A1 => n14252, A2 => n14253, A3 => n14254, A4 => 
                           n14255, ZN => n14251);
   U8730 : NOR2_X1 port map( A1 => n14251, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N164);
   U8849 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_31_25_port,
                           A2 => n17154, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_25_port, B2 => 
                           n17683, ZN => n14368);
   U8848 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_29_25_port,
                           A2 => n17684, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_25_port, B2 => 
                           n17685, ZN => n14369);
   U8847 : AOI222_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_4_25_port,
                           A2 => n17686, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_25_port, B2 => 
                           n17153, C1 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_25_port, C2 => 
                           n17687, ZN => n14370);
   U8846 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_27_25_port,
                           A2 => n17688, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_25_port, B2 => 
                           n17689, ZN => n14364);
   U8845 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_23_25_port,
                           A2 => n17690, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_25_port, B2 => 
                           n17691, ZN => n14365);
   U8844 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_21_25_port,
                           A2 => n17692, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_25_port, B2 => 
                           n17693, ZN => n14366);
   U8843 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_19_25_port,
                           A2 => n17694, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_25_port, B2 => 
                           n17695, ZN => n14367);
   U8842 : NAND4_X1 port map( A1 => n14364, A2 => n14365, A3 => n14366, A4 => 
                           n14367, ZN => n14353);
   U8841 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_17_25_port,
                           A2 => n17696, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_25_port, B2 => 
                           n17697, ZN => n14360);
   U8840 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_12_25_port,
                           A2 => n17698, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_25_port, B2 => 
                           n17357, ZN => n14361);
   U8839 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_8_25_port, 
                           A2 => n17417, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_25_port, B2 => 
                           n17152, ZN => n14362);
   U8838 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_9_25_port, 
                           A2 => n17351, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_25_port, B2 => 
                           n17699, ZN => n14363);
   U8837 : NAND4_X1 port map( A1 => n14360, A2 => n14361, A3 => n14362, A4 => 
                           n14363, ZN => n14354);
   U8836 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_11_25_port,
                           A2 => n17151, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_25_port, B2 => 
                           n17413, ZN => n14356);
   U8835 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_14_25_port,
                           A2 => n17700, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_25_port, B2 => 
                           n17414, ZN => n14357);
   U8834 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_2_25_port, 
                           A2 => n17353, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_25_port, B2 => 
                           n17415, ZN => n14358);
   U8833 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_6_25_port, 
                           A2 => n17354, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_25_port, B2 => 
                           n17416, ZN => n14359);
   U8832 : NAND4_X1 port map( A1 => n14356, A2 => n14357, A3 => n14358, A4 => 
                           n14359, ZN => n14355);
   U8831 : NOR4_X1 port map( A1 => n14352, A2 => n14353, A3 => n14354, A4 => 
                           n14355, ZN => n14351);
   U8830 : NOR2_X1 port map( A1 => n14351, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N159);
   U9289 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_31_3_port, 
                           A2 => n17154, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_30_3_port, B2 => 
                           n17683, ZN => n14808);
   U9288 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_29_3_port, 
                           A2 => n14247, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_28_3_port, B2 => 
                           n17685, ZN => n14809);
   U9287 : AOI222_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_4_3_port, 
                           A2 => n17686, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_25_3_port, B2 => 
                           n17153, C1 => 
                           pipeline_RegFile_DEC_WB_RegBank_24_3_port, C2 => 
                           n17687, ZN => n14810);
   U9286 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_27_3_port, 
                           A2 => n17688, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_26_3_port, B2 => 
                           n17689, ZN => n14804);
   U9285 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_23_3_port, 
                           A2 => n17690, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_22_3_port, B2 => 
                           n17691, ZN => n14805);
   U9284 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_21_3_port, 
                           A2 => n17692, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_20_3_port, B2 => 
                           n17693, ZN => n14806);
   U9283 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_19_3_port, 
                           A2 => n14233, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_18_3_port, B2 => 
                           n17695, ZN => n14807);
   U9282 : NAND4_X1 port map( A1 => n14804, A2 => n14805, A3 => n14806, A4 => 
                           n14807, ZN => n14793);
   U9281 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_17_3_port, 
                           A2 => n17696, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_16_3_port, B2 => 
                           n17697, ZN => n14800);
   U9280 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_12_3_port, 
                           A2 => n17698, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_13_3_port, B2 => 
                           n17357, ZN => n14801);
   U9279 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_8_3_port, 
                           A2 => n17417, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_15_3_port, B2 => 
                           n17152, ZN => n14802);
   U9278 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_9_3_port, 
                           A2 => n17351, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_10_3_port, B2 => 
                           n17699, ZN => n14803);
   U9277 : NAND4_X1 port map( A1 => n14800, A2 => n14801, A3 => n14802, A4 => 
                           n14803, ZN => n14794);
   U9276 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_11_3_port, 
                           A2 => n17151, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_3_3_port, B2 => 
                           n17413, ZN => n14796);
   U9275 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_14_3_port, 
                           A2 => n17700, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_5_3_port, B2 => 
                           n17414, ZN => n14797);
   U9274 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_2_3_port, 
                           A2 => n17353, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_7_3_port, B2 => 
                           n17415, ZN => n14798);
   U9273 : AOI22_X1 port map( A1 => pipeline_RegFile_DEC_WB_RegBank_6_3_port, 
                           A2 => n17354, B1 => 
                           pipeline_RegFile_DEC_WB_RegBank_1_3_port, B2 => 
                           n17416, ZN => n14799);
   U9272 : NAND4_X1 port map( A1 => n14796, A2 => n14797, A3 => n14798, A4 => 
                           n14799, ZN => n14795);
   U9271 : NOR4_X1 port map( A1 => n14792, A2 => n14793, A3 => n14794, A4 => 
                           n14795, ZN => n14791);
   U9270 : NOR2_X1 port map( A1 => n14791, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N137);
   U9420 : OAI22_X1 port map( A1 => n14913, A2 => n17075, B1 => n17109, B2 => 
                           n17461, ZN => pipeline_IDEX_Stage_N118);
   U9402 : OAI22_X1 port map( A1 => n14895, A2 => n17075, B1 => n17682, B2 => 
                           n17451, ZN => pipeline_IDEX_Stage_N127);
   U9452 : OAI22_X1 port map( A1 => n14945, A2 => n17075, B1 => n17109, B2 => 
                           n17450, ZN => pipeline_IDEX_Stage_N102);
   U9442 : OAI22_X1 port map( A1 => n14935, A2 => n17075, B1 => n17109, B2 => 
                           n17454, ZN => pipeline_IDEX_Stage_N107);
   U9414 : OAI22_X1 port map( A1 => n14907, A2 => n17075, B1 => n17109, B2 => 
                           n17438, ZN => pipeline_IDEX_Stage_N121);
   U9390 : OAI22_X1 port map( A1 => n14883, A2 => n17075, B1 => n17109, B2 => 
                           n17527, ZN => pipeline_IDEX_Stage_N133);
   U8698 : NOR2_X1 port map( A1 => n17350, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N171);
   U8668 : NOR2_X1 port map( A1 => n17349, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N206);
   U8686 : NOR2_X1 port map( A1 => n17433, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N177);
   U8696 : NOR2_X1 port map( A1 => n17361, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N172);
   U8702 : NOR2_X1 port map( A1 => n17410, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N169);
   U8706 : NOR2_X1 port map( A1 => n17406, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N167);
   U8684 : NOR2_X1 port map( A1 => n17444, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N178);
   U8674 : NOR2_X1 port map( A1 => n17383, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N200);
   U8694 : NOR2_X1 port map( A1 => n17437, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N173);
   U8669 : NOR2_X1 port map( A1 => n17408, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N205);
   U8672 : NOR2_X1 port map( A1 => n17328, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N202);
   U8673 : NOR2_X1 port map( A1 => n17384, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N201);
   U8671 : NOR2_X1 port map( A1 => n17316, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N203);
   U9394 : OAI22_X1 port map( A1 => n14887, A2 => n17075, B1 => n17109, B2 => 
                           n17452, ZN => pipeline_IDEX_Stage_N131);
   U9422 : OAI22_X1 port map( A1 => n14915, A2 => n17075, B1 => n17109, B2 => 
                           n17453, ZN => pipeline_IDEX_Stage_N117);
   U9424 : OAI22_X1 port map( A1 => n14917, A2 => n17075, B1 => n17682, B2 => 
                           n17460, ZN => pipeline_IDEX_Stage_N116);
   U8690 : NOR2_X1 port map( A1 => n17432, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N175);
   U8675 : NOR2_X1 port map( A1 => n17317, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N199);
   U8708 : NOR2_X1 port map( A1 => n17076, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N166);
   U8682 : NOR2_X1 port map( A1 => n17434, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N179);
   U8692 : NOR2_X1 port map( A1 => n17428, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N174);
   U8680 : NOR2_X1 port map( A1 => n17445, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N180);
   U8700 : NOR2_X1 port map( A1 => n17412, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N170);
   U8670 : NOR2_X1 port map( A1 => n17329, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N204);
   U8667 : NOR2_X1 port map( A1 => n17407, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N207);
   U8676 : NOR2_X1 port map( A1 => n17315, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N198);
   U8688 : NOR2_X1 port map( A1 => n17440, A2 => n17075, ZN => 
                           pipeline_IDEX_Stage_N176);
   U8594 : AOI22_X1 port map( A1 => pipeline_Alu_Out_Addr_to_mem_1_port, A2 => 
                           n17370, B1 => n14135, B2 => data_from_dram_1_port, 
                           ZN => n14165);
   U8596 : AOI22_X1 port map( A1 => pipeline_Alu_Out_Addr_to_mem_0_port, A2 => 
                           n17370, B1 => n14135, B2 => data_from_dram_0_port, 
                           ZN => n14166);
   U8566 : AOI22_X1 port map( A1 => pipeline_Alu_Out_Addr_to_mem_15_port, A2 =>
                           n14134, B1 => n14135, B2 => data_from_dram_15_port, 
                           ZN => n14151);
   U8570 : AOI22_X1 port map( A1 => pipeline_Alu_Out_Addr_to_mem_13_port, A2 =>
                           n14134, B1 => n14135, B2 => data_from_dram_13_port, 
                           ZN => n14153);
   U8548 : AOI22_X1 port map( A1 => pipeline_Alu_Out_Addr_to_mem_24_port, A2 =>
                           n17370, B1 => n14135, B2 => data_from_dram_24_port, 
                           ZN => n14142);
   U8584 : AOI22_X1 port map( A1 => pipeline_Alu_Out_Addr_to_mem_6_port, A2 => 
                           n17370, B1 => n14135, B2 => data_from_dram_6_port, 
                           ZN => n14160);
   U8540 : AOI22_X1 port map( A1 => pipeline_Alu_Out_Addr_to_mem_28_port, A2 =>
                           n17370, B1 => n14135, B2 => data_from_dram_28_port, 
                           ZN => n14138);
   U8572 : AOI22_X1 port map( A1 => pipeline_Alu_Out_Addr_to_mem_12_port, A2 =>
                           n14134, B1 => n14135, B2 => data_from_dram_12_port, 
                           ZN => n14154);
   U8534 : AOI22_X1 port map( A1 => pipeline_Alu_Out_Addr_to_mem_31_port, A2 =>
                           n14134, B1 => n14135, B2 => data_from_dram_31_port, 
                           ZN => n14133);
   U8546 : AOI22_X1 port map( A1 => pipeline_Alu_Out_Addr_to_mem_25_port, A2 =>
                           n17370, B1 => n14135, B2 => data_from_dram_25_port, 
                           ZN => n14141);
   U8550 : AOI22_X1 port map( A1 => pipeline_Alu_Out_Addr_to_mem_23_port, A2 =>
                           n17370, B1 => n14135, B2 => data_from_dram_23_port, 
                           ZN => n14143);
   U8588 : AOI22_X1 port map( A1 => pipeline_Alu_Out_Addr_to_mem_4_port, A2 => 
                           n17370, B1 => n14135, B2 => data_from_dram_4_port, 
                           ZN => n14162);
   U8590 : AOI22_X1 port map( A1 => pipeline_Alu_Out_Addr_to_mem_3_port, A2 => 
                           n17370, B1 => n14135, B2 => data_from_dram_3_port, 
                           ZN => n14163);
   U8580 : AOI22_X1 port map( A1 => pipeline_Alu_Out_Addr_to_mem_8_port, A2 => 
                           n17370, B1 => n14135, B2 => data_from_dram_8_port, 
                           ZN => n14158);
   U8582 : AOI22_X1 port map( A1 => pipeline_Alu_Out_Addr_to_mem_7_port, A2 => 
                           n17370, B1 => n14135, B2 => data_from_dram_7_port, 
                           ZN => n14159);
   U8552 : AOI22_X1 port map( A1 => pipeline_Alu_Out_Addr_to_mem_22_port, A2 =>
                           n17370, B1 => n14135, B2 => data_from_dram_22_port, 
                           ZN => n14144);
   U8592 : AOI22_X1 port map( A1 => pipeline_Alu_Out_Addr_to_mem_2_port, A2 => 
                           n17370, B1 => n14135, B2 => data_from_dram_2_port, 
                           ZN => n14164);
   U8578 : AOI22_X1 port map( A1 => pipeline_Alu_Out_Addr_to_mem_9_port, A2 => 
                           n14134, B1 => n14135, B2 => data_from_dram_9_port, 
                           ZN => n14157);
   U8554 : AOI22_X1 port map( A1 => pipeline_Alu_Out_Addr_to_mem_21_port, A2 =>
                           n14134, B1 => n14135, B2 => data_from_dram_21_port, 
                           ZN => n14145);
   U8574 : AOI22_X1 port map( A1 => pipeline_Alu_Out_Addr_to_mem_11_port, A2 =>
                           n14134, B1 => n14135, B2 => data_from_dram_11_port, 
                           ZN => n14155);
   U8560 : AOI22_X1 port map( A1 => pipeline_Alu_Out_Addr_to_mem_18_port, A2 =>
                           n14134, B1 => n14135, B2 => data_from_dram_18_port, 
                           ZN => n14148);
   U8556 : AOI22_X1 port map( A1 => pipeline_Alu_Out_Addr_to_mem_20_port, A2 =>
                           n14134, B1 => n14135, B2 => data_from_dram_20_port, 
                           ZN => n14146);
   U8536 : AOI22_X1 port map( A1 => pipeline_Alu_Out_Addr_to_mem_30_port, A2 =>
                           n17370, B1 => n14135, B2 => data_from_dram_30_port, 
                           ZN => n14136);
   U8538 : AOI22_X1 port map( A1 => pipeline_Alu_Out_Addr_to_mem_29_port, A2 =>
                           n17370, B1 => n14135, B2 => data_from_dram_29_port, 
                           ZN => n14137);
   U8542 : AOI22_X1 port map( A1 => pipeline_Alu_Out_Addr_to_mem_27_port, A2 =>
                           n17370, B1 => n14135, B2 => data_from_dram_27_port, 
                           ZN => n14139);
   U8558 : AOI22_X1 port map( A1 => pipeline_Alu_Out_Addr_to_mem_19_port, A2 =>
                           n14134, B1 => n14135, B2 => data_from_dram_19_port, 
                           ZN => n14147);
   U8544 : AOI22_X1 port map( A1 => pipeline_Alu_Out_Addr_to_mem_26_port, A2 =>
                           n17370, B1 => n14135, B2 => data_from_dram_26_port, 
                           ZN => n14140);
   U8568 : AOI22_X1 port map( A1 => pipeline_Alu_Out_Addr_to_mem_14_port, A2 =>
                           n14134, B1 => n14135, B2 => data_from_dram_14_port, 
                           ZN => n14152);
   U8586 : AOI22_X1 port map( A1 => pipeline_Alu_Out_Addr_to_mem_5_port, A2 => 
                           n17370, B1 => n14135, B2 => data_from_dram_5_port, 
                           ZN => n14161);
   U8562 : AOI22_X1 port map( A1 => pipeline_Alu_Out_Addr_to_mem_17_port, A2 =>
                           n14134, B1 => n14135, B2 => data_from_dram_17_port, 
                           ZN => n14149);
   U8564 : AOI22_X1 port map( A1 => pipeline_Alu_Out_Addr_to_mem_16_port, A2 =>
                           n14134, B1 => n14135, B2 => data_from_dram_16_port, 
                           ZN => n14150);
   U8576 : AOI22_X1 port map( A1 => pipeline_Alu_Out_Addr_to_mem_10_port, A2 =>
                           n14134, B1 => n14135, B2 => data_from_dram_10_port, 
                           ZN => n14156);
   U8608 : NAND2_X1 port map( A1 => n17703, A2 => n14007, ZN => n13988);
   U8607 : NOR2_X1 port map( A1 => n14168, A2 => n13988, ZN => 
                           pipeline_IDEX_Stage_N92);
   U8611 : NOR2_X1 port map( A1 => n17382, A2 => n14169, ZN => n14123);
   U8609 : NOR2_X1 port map( A1 => n14168, A2 => n13981, ZN => 
                           pipeline_IDEX_Stage_N91);
   U8663 : AOI21_X1 port map( B1 => n14025, B2 => n17349, A => n14168, ZN => 
                           pipeline_IDEX_Stage_N211);
   U8704 : AOI21_X1 port map( B1 => n14025, B2 => n17404, A => n14168, ZN => 
                           pipeline_IDEX_Stage_N168);
   U8664 : AOI21_X1 port map( B1 => n14025, B2 => n17408, A => n14168, ZN => 
                           pipeline_IDEX_Stage_N210);
   U8659 : AOI21_X1 port map( B1 => n14025, B2 => n17434, A => n14168, ZN => 
                           pipeline_IDEX_Stage_N215);
   U8657 : AOI21_X1 port map( B1 => n14025, B2 => n17431, A => n14168, ZN => 
                           pipeline_IDEX_Stage_N217);
   U8658 : AOI21_X1 port map( B1 => n14025, B2 => n17445, A => n14168, ZN => 
                           pipeline_IDEX_Stage_N216);
   U8662 : AOI21_X1 port map( B1 => n14025, B2 => n17407, A => n14168, ZN => 
                           pipeline_IDEX_Stage_N212);
   U8666 : AOI21_X1 port map( B1 => n14025, B2 => n17316, A => n14168, ZN => 
                           pipeline_IDEX_Stage_N208);
   U8665 : AOI21_X1 port map( B1 => n14025, B2 => n17329, A => n14168, ZN => 
                           pipeline_IDEX_Stage_N209);
   U8660 : AOI21_X1 port map( B1 => n14025, B2 => n17444, A => n14168, ZN => 
                           pipeline_IDEX_Stage_N214);
   U8661 : AOI21_X1 port map( B1 => n14025, B2 => n17433, A => n14168, ZN => 
                           pipeline_IDEX_Stage_N213);
   U9474 : NOR3_X1 port map( A1 => n14982, A2 => n17447, A3 => n14129, ZN => 
                           pipeline_EXMEM_stage_N76);
   U8528 : NOR2_X1 port map( A1 => n17393, A2 => n14129, ZN => 
                           pipeline_MEMWB_Stage_N47);
   U8531 : NOR2_X1 port map( A1 => n17645, A2 => n14129, ZN => 
                           pipeline_MEMWB_Stage_N44);
   U8530 : NOR2_X1 port map( A1 => n17646, A2 => n14129, ZN => 
                           pipeline_MEMWB_Stage_N45);
   U9476 : NOR2_X1 port map( A1 => Rst, A2 => n14101, ZN => 
                           pipeline_EXMEM_stage_N75);
   U9483 : AOI22_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_7_port, A2
                           => n13931, B1 => n13926, B2 => n17430, ZN => n14117)
                           ;
   U9482 : NOR2_X1 port map( A1 => Rst, A2 => n14117, ZN => 
                           pipeline_EXMEM_stage_N72);
   U9485 : AOI22_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_7_port, A2
                           => n13930, B1 => n13925, B2 => n17430, ZN => n14116)
                           ;
   U9484 : NOR2_X1 port map( A1 => Rst, A2 => n14116, ZN => 
                           pipeline_EXMEM_stage_N71);
   U10044 : OAI21_X1 port map( B1 => n15646, B2 => n17371, A => n17703, ZN => 
                           n3925);
   U10042 : OAI21_X1 port map( B1 => n15646, B2 => n17372, A => n17703, ZN => 
                           n3926);
   U10022 : OAI21_X1 port map( B1 => n15646, B2 => n17478, A => n17702, ZN => 
                           n3936);
   U10038 : OAI21_X1 port map( B1 => n15646, B2 => n17472, A => n17702, ZN => 
                           n3928);
   U10016 : OAI21_X1 port map( B1 => n15646, B2 => n17481, A => n17702, ZN => 
                           n3939);
   U10018 : OAI21_X1 port map( B1 => n15646, B2 => n17480, A => n17702, ZN => 
                           n3938);
   U10020 : OAI21_X1 port map( B1 => n15646, B2 => n17479, A => n17702, ZN => 
                           n3937);
   U10026 : OAI21_X1 port map( B1 => n15646, B2 => n17477, A => n17702, ZN => 
                           n3934);
   U10028 : OAI21_X1 port map( B1 => n15646, B2 => n17476, A => n17702, ZN => 
                           n3933);
   U10024 : OAI21_X1 port map( B1 => n15646, B2 => n17375, A => n17701, ZN => 
                           n3935);
   U10004 : OAI21_X1 port map( B1 => n15646, B2 => n17378, A => n17701, ZN => 
                           n3945);
   U10002 : OAI21_X1 port map( B1 => n15646, B2 => n17485, A => n17701, ZN => 
                           n3946);
   U10000 : OAI21_X1 port map( B1 => n15646, B2 => n17486, A => n17701, ZN => 
                           n3947);
   U9998 : OAI21_X1 port map( B1 => n15646, B2 => n17487, A => n17701, ZN => 
                           n3948);
   U9996 : OAI21_X1 port map( B1 => n15646, B2 => n17488, A => n17701, ZN => 
                           n3949);
   U9994 : OAI21_X1 port map( B1 => n15646, B2 => n17489, A => n17701, ZN => 
                           n3950);
   U9992 : OAI21_X1 port map( B1 => n15646, B2 => n17490, A => n17701, ZN => 
                           n3951);
   U9990 : OAI21_X1 port map( B1 => n15646, B2 => n17491, A => n17701, ZN => 
                           n3952);
   U10014 : OAI21_X1 port map( B1 => n15646, B2 => n17376, A => n17702, ZN => 
                           n3940);
   U10012 : OAI21_X1 port map( B1 => n15646, B2 => n17377, A => n17701, ZN => 
                           n3941);
   U10010 : OAI21_X1 port map( B1 => n15646, B2 => n17482, A => n17701, ZN => 
                           n3942);
   U10008 : OAI21_X1 port map( B1 => n15646, B2 => n17483, A => n17701, ZN => 
                           n3943);
   U10006 : OAI21_X1 port map( B1 => n15646, B2 => n17484, A => n17701, ZN => 
                           n3944);
   U10030 : OAI21_X1 port map( B1 => n15646, B2 => n17475, A => n17702, ZN => 
                           n3932);
   U10032 : OAI21_X1 port map( B1 => n15646, B2 => n17474, A => n17702, ZN => 
                           n3931);
   U10034 : OAI21_X1 port map( B1 => n15646, B2 => n17473, A => n17702, ZN => 
                           n3930);
   U10036 : OAI21_X1 port map( B1 => n15646, B2 => n17374, A => n17702, ZN => 
                           n3929);
   U10040 : OAI21_X1 port map( B1 => n15646, B2 => n17373, A => n17702, ZN => 
                           n3927);
   U9481 : AOI22_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_7_port, A2
                           => n13932, B1 => n13927, B2 => n17430, ZN => n14113)
                           ;
   U9480 : NOR2_X1 port map( A1 => Rst, A2 => n14113, ZN => 
                           pipeline_EXMEM_stage_N73);
   U9479 : AOI22_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_7_port, A2
                           => n13933, B1 => n13928, B2 => n17430, ZN => n14100)
                           ;
   U9478 : NOR2_X1 port map( A1 => Rst, A2 => n14100, ZN => 
                           pipeline_EXMEM_stage_N74);
   U9984 : OAI21_X1 port map( B1 => n15646, B2 => n17494, A => n17701, ZN => 
                           n3955);
   U9982 : OAI21_X1 port map( B1 => n15646, B2 => n17379, A => n17702, ZN => 
                           n3956);
   U9986 : OAI21_X1 port map( B1 => n15646, B2 => n17493, A => n17702, ZN => 
                           n3954);
   U9988 : OAI21_X1 port map( B1 => n15646, B2 => n17492, A => n17705, ZN => 
                           n3953);
   U9563 : NOR2_X1 port map( A1 => Rst, A2 => n17447, ZN => 
                           pipeline_EXMEM_stage_N5);
   U9585 : NOR2_X1 port map( A1 => Rst, A2 => n17449, ZN => 
                           pipeline_EXMEM_stage_N4);
   U11058 : OAI21_X1 port map( B1 => n15001, B2 => n16598, A => 
                           pipeline_EXE_controls_in_EXEcute_5_port, ZN => 
                           n16599);
   U11057 : AOI211_X1 port map( C1 => n15001, C2 => n16598, A => 
                           pipeline_EXE_controls_in_EXEcute_6_port, B => n16599
                           , ZN => exception);
   U11949 : NOR2_X1 port map( A1 => n17000, A2 => n16597, ZN => DataMem_N1671);
   U11894 : NOR2_X1 port map( A1 => n17000, A2 => n16596, ZN => DataMem_N1735);
   U11859 : NOR2_X1 port map( A1 => n17000, A2 => n16595, ZN => DataMem_N1799);
   U11599 : AOI22_X1 port map( A1 => n16823, A2 => DataMem_Mem_7_11_port, B1 =>
                           n16824, B2 => DataMem_Mem_6_11_port, ZN => n16921);
   U11769 : NAND2_X1 port map( A1 => addr_to_dataRam_4_port, A2 => 
                           addr_to_dataRam_2_port, ZN => n17014);
   U11598 : AOI22_X1 port map( A1 => n16821, A2 => DataMem_Mem_5_11_port, B1 =>
                           n16822, B2 => DataMem_Mem_4_11_port, ZN => n16922);
   U11838 : NAND2_X1 port map( A1 => addr_to_dataRam_2_port, A2 => 
                           addr_to_dataRam_3_port, ZN => n17016);
   U11872 : NOR3_X1 port map( A1 => addr_to_dataRam_4_port, A2 => 
                           addr_to_dataRam_2_port, A3 => n17015, ZN => n16820);
   U11597 : AOI22_X1 port map( A1 => n17122, A2 => DataMem_Mem_3_11_port, B1 =>
                           n17653, B2 => DataMem_Mem_2_11_port, ZN => n16923);
   U11596 : AOI22_X1 port map( A1 => n17124, A2 => DataMem_Mem_1_11_port, B1 =>
                           n17125, B2 => DataMem_Mem_0_11_port, ZN => n16924);
   U11594 : NOR2_X1 port map( A1 => n17155, A2 => n16920, ZN => DataMem_N2194);
   U11687 : NOR2_X1 port map( A1 => n17001, A2 => n16590, ZN => DataMem_N2117);
   U11721 : NOR2_X1 port map( A1 => n17001, A2 => n16591, ZN => DataMem_N2053);
   U11756 : NOR2_X1 port map( A1 => n17001, A2 => n16592, ZN => DataMem_N1989);
   U11791 : NOR2_X1 port map( A1 => n17001, A2 => n16593, ZN => DataMem_N1925);
   U11825 : NOR2_X1 port map( A1 => n17001, A2 => n16594, ZN => DataMem_N1861);
   U11860 : NOR2_X1 port map( A1 => n17001, A2 => n16595, ZN => DataMem_N1797);
   U11895 : NOR2_X1 port map( A1 => n17001, A2 => n16596, ZN => DataMem_N1733);
   U11947 : NOR2_X1 port map( A1 => n16999, A2 => n17650, ZN => DataMem_N1673);
   U11593 : AOI22_X1 port map( A1 => n16823, A2 => DataMem_Mem_7_12_port, B1 =>
                           n16824, B2 => DataMem_Mem_6_12_port, ZN => n16916);
   U11592 : AOI22_X1 port map( A1 => n16821, A2 => DataMem_Mem_5_12_port, B1 =>
                           n16822, B2 => DataMem_Mem_4_12_port, ZN => n16917);
   U11591 : AOI22_X1 port map( A1 => n17122, A2 => DataMem_Mem_3_12_port, B1 =>
                           n17653, B2 => DataMem_Mem_2_12_port, ZN => n16918);
   U11590 : AOI22_X1 port map( A1 => n17124, A2 => DataMem_Mem_1_12_port, B1 =>
                           n17125, B2 => DataMem_Mem_0_12_port, ZN => n16919);
   U11588 : NOR2_X1 port map( A1 => n17155, A2 => n16915, ZN => DataMem_N2197);
   U11695 : NOR2_X1 port map( A1 => n17009, A2 => n17661, ZN => DataMem_N2101);
   U11729 : NOR2_X1 port map( A1 => n17009, A2 => n17658, ZN => DataMem_N2037);
   U11764 : NOR2_X1 port map( A1 => n17009, A2 => n17657, ZN => DataMem_N1973);
   U11799 : NOR2_X1 port map( A1 => n17009, A2 => n17656, ZN => DataMem_N1909);
   U11833 : NOR2_X1 port map( A1 => n17009, A2 => n17655, ZN => DataMem_N1845);
   U11868 : NOR2_X1 port map( A1 => n17009, A2 => n17654, ZN => DataMem_N1781);
   U11903 : NOR2_X1 port map( A1 => n17009, A2 => n17651, ZN => DataMem_N1717);
   U11967 : NOR2_X1 port map( A1 => n17009, A2 => n17650, ZN => DataMem_N1653);
   U11940 : AOI22_X1 port map( A1 => pipeline_Forward_sw1_mux, A2 => 
                           pipeline_data_to_RF_from_WB_16_port, B1 => n13803, 
                           B2 => n17380, ZN => n16995);
   U11854 : NOR2_X1 port map( A1 => n16995, A2 => n17654, ZN => DataMem_N1809);
   U11653 : AOI22_X1 port map( A1 => n17659, A2 => DataMem_Mem_7_2_port, B1 => 
                           n17530, B2 => DataMem_Mem_6_2_port, ZN => n16966);
   U11652 : AOI22_X1 port map( A1 => n17531, A2 => DataMem_Mem_5_2_port, B1 => 
                           n16822, B2 => DataMem_Mem_4_2_port, ZN => n16967);
   U11651 : AOI22_X1 port map( A1 => n17122, A2 => DataMem_Mem_3_2_port, B1 => 
                           n17653, B2 => DataMem_Mem_2_2_port, ZN => n16968);
   U11650 : AOI22_X1 port map( A1 => n17124, A2 => DataMem_Mem_1_2_port, B1 => 
                           n17125, B2 => DataMem_Mem_0_2_port, ZN => n16969);
   U11648 : NOR2_X1 port map( A1 => n17155, A2 => n16965, ZN => DataMem_N2167);
   U11694 : NOR2_X1 port map( A1 => n17008, A2 => n17661, ZN => DataMem_N2103);
   U11728 : NOR2_X1 port map( A1 => n17008, A2 => n17658, ZN => DataMem_N2039);
   U11763 : NOR2_X1 port map( A1 => n17008, A2 => n17657, ZN => DataMem_N1975);
   U11798 : NOR2_X1 port map( A1 => n17008, A2 => n17656, ZN => DataMem_N1911);
   U11832 : NOR2_X1 port map( A1 => n17008, A2 => n17655, ZN => DataMem_N1847);
   U11867 : NOR2_X1 port map( A1 => n17008, A2 => n17654, ZN => DataMem_N1783);
   U11902 : NOR2_X1 port map( A1 => n17008, A2 => n17651, ZN => DataMem_N1719);
   U11965 : NOR2_X1 port map( A1 => n17008, A2 => n17650, ZN => DataMem_N1655);
   U11647 : AOI22_X1 port map( A1 => n17660, A2 => DataMem_Mem_7_3_port, B1 => 
                           n17530, B2 => DataMem_Mem_6_3_port, ZN => n16961);
   U11646 : AOI22_X1 port map( A1 => n17531, A2 => DataMem_Mem_5_3_port, B1 => 
                           n16822, B2 => DataMem_Mem_4_3_port, ZN => n16962);
   U11645 : AOI22_X1 port map( A1 => n17122, A2 => DataMem_Mem_3_3_port, B1 => 
                           n17653, B2 => DataMem_Mem_2_3_port, ZN => n16963);
   U11644 : AOI22_X1 port map( A1 => n17124, A2 => DataMem_Mem_1_3_port, B1 => 
                           n17125, B2 => DataMem_Mem_0_3_port, ZN => n16964);
   U11642 : NOR2_X1 port map( A1 => n17155, A2 => n16960, ZN => DataMem_N2170);
   U11681 : NOR2_X1 port map( A1 => n16995, A2 => n17661, ZN => DataMem_N2129);
   U11715 : NOR2_X1 port map( A1 => n16995, A2 => n17658, ZN => DataMem_N2065);
   U11750 : NOR2_X1 port map( A1 => n16995, A2 => n17657, ZN => DataMem_N2001);
   U11785 : NOR2_X1 port map( A1 => n16995, A2 => n17656, ZN => DataMem_N1937);
   U11819 : NOR2_X1 port map( A1 => n16995, A2 => n17655, ZN => DataMem_N1873);
   U11685 : NOR2_X1 port map( A1 => n16999, A2 => n17661, ZN => DataMem_N2121);
   U11719 : NOR2_X1 port map( A1 => n16999, A2 => n17658, ZN => DataMem_N2057);
   U11754 : NOR2_X1 port map( A1 => n16999, A2 => n17657, ZN => DataMem_N1993);
   U11789 : NOR2_X1 port map( A1 => n16999, A2 => n17656, ZN => DataMem_N1929);
   U11823 : NOR2_X1 port map( A1 => n16999, A2 => n17655, ZN => DataMem_N1865);
   U11858 : NOR2_X1 port map( A1 => n16999, A2 => n17654, ZN => DataMem_N1801);
   U11893 : NOR2_X1 port map( A1 => n16999, A2 => n17651, ZN => DataMem_N1737);
   U11696 : NOR2_X1 port map( A1 => n17010, A2 => n17661, ZN => DataMem_N2099);
   U11730 : NOR2_X1 port map( A1 => n17010, A2 => n17658, ZN => DataMem_N2035);
   U11765 : NOR2_X1 port map( A1 => n17010, A2 => n17657, ZN => DataMem_N1971);
   U11800 : NOR2_X1 port map( A1 => n17010, A2 => n17656, ZN => DataMem_N1907);
   U11834 : NOR2_X1 port map( A1 => n17010, A2 => n17655, ZN => DataMem_N1843);
   U11869 : NOR2_X1 port map( A1 => n17010, A2 => n17654, ZN => DataMem_N1779);
   U11904 : NOR2_X1 port map( A1 => n17010, A2 => n17651, ZN => DataMem_N1715);
   U11759 : NOR2_X1 port map( A1 => n17004, A2 => n17657, ZN => DataMem_N1983);
   U11693 : NOR2_X1 port map( A1 => n17007, A2 => n17661, ZN => DataMem_N2105);
   U11727 : NOR2_X1 port map( A1 => n17007, A2 => n17658, ZN => DataMem_N2041);
   U11762 : NOR2_X1 port map( A1 => n17007, A2 => n17657, ZN => DataMem_N1977);
   U11797 : NOR2_X1 port map( A1 => n17007, A2 => n17656, ZN => DataMem_N1913);
   U11831 : NOR2_X1 port map( A1 => n17007, A2 => n17655, ZN => DataMem_N1849);
   U11866 : NOR2_X1 port map( A1 => n17007, A2 => n17654, ZN => DataMem_N1785);
   U11901 : NOR2_X1 port map( A1 => n17007, A2 => n17651, ZN => DataMem_N1721);
   U11963 : NOR2_X1 port map( A1 => n17007, A2 => n17650, ZN => DataMem_N1657);
   U11641 : AOI22_X1 port map( A1 => n17660, A2 => DataMem_Mem_7_4_port, B1 => 
                           n17530, B2 => DataMem_Mem_6_4_port, ZN => n16956);
   U11640 : AOI22_X1 port map( A1 => n17531, A2 => DataMem_Mem_5_4_port, B1 => 
                           n16822, B2 => DataMem_Mem_4_4_port, ZN => n16957);
   U11639 : AOI22_X1 port map( A1 => n17122, A2 => DataMem_Mem_3_4_port, B1 => 
                           n17652, B2 => DataMem_Mem_2_4_port, ZN => n16958);
   U11638 : AOI22_X1 port map( A1 => n17124, A2 => DataMem_Mem_1_4_port, B1 => 
                           n17125, B2 => DataMem_Mem_0_4_port, ZN => n16959);
   U11636 : NOR2_X1 port map( A1 => n17155, A2 => n16955, ZN => DataMem_N2173);
   U11605 : AOI22_X1 port map( A1 => n16823, A2 => DataMem_Mem_7_10_port, B1 =>
                           n16824, B2 => DataMem_Mem_6_10_port, ZN => n16926);
   U11604 : AOI22_X1 port map( A1 => n16821, A2 => DataMem_Mem_5_10_port, B1 =>
                           n16822, B2 => DataMem_Mem_4_10_port, ZN => n16927);
   U11603 : AOI22_X1 port map( A1 => n17122, A2 => DataMem_Mem_3_10_port, B1 =>
                           n17653, B2 => DataMem_Mem_2_10_port, ZN => n16928);
   U11602 : AOI22_X1 port map( A1 => n17124, A2 => DataMem_Mem_1_10_port, B1 =>
                           n17125, B2 => DataMem_Mem_0_10_port, ZN => n16929);
   U11600 : NOR2_X1 port map( A1 => n17155, A2 => n16925, ZN => DataMem_N2191);
   U11951 : NOR2_X1 port map( A1 => n17001, A2 => n16597, ZN => DataMem_N1669);
   U11899 : NOR2_X1 port map( A1 => n17005, A2 => n17651, ZN => DataMem_N1725);
   U11864 : NOR2_X1 port map( A1 => n17005, A2 => n17654, ZN => DataMem_N1789);
   U11829 : NOR2_X1 port map( A1 => n17005, A2 => n17655, ZN => DataMem_N1853);
   U11795 : NOR2_X1 port map( A1 => n17005, A2 => n17656, ZN => DataMem_N1917);
   U11760 : NOR2_X1 port map( A1 => n17005, A2 => n17657, ZN => DataMem_N1981);
   U11725 : NOR2_X1 port map( A1 => n17005, A2 => n17658, ZN => DataMem_N2045);
   U11691 : NOR2_X1 port map( A1 => n17005, A2 => n17661, ZN => DataMem_N2109);
   U11623 : AOI22_X1 port map( A1 => n16823, A2 => DataMem_Mem_7_7_port, B1 => 
                           n16824, B2 => DataMem_Mem_6_7_port, ZN => n16941);
   U11622 : AOI22_X1 port map( A1 => n17531, A2 => DataMem_Mem_5_7_port, B1 => 
                           n16822, B2 => DataMem_Mem_4_7_port, ZN => n16942);
   U11621 : AOI22_X1 port map( A1 => n16819, A2 => DataMem_Mem_3_7_port, B1 => 
                           n17653, B2 => DataMem_Mem_2_7_port, ZN => n16943);
   U11620 : AOI22_X1 port map( A1 => n17124, A2 => DataMem_Mem_1_7_port, B1 => 
                           n17125, B2 => DataMem_Mem_0_7_port, ZN => n16944);
   U11618 : NOR2_X1 port map( A1 => n17155, A2 => n16940, ZN => DataMem_N2182);
   U11957 : NOR2_X1 port map( A1 => n17004, A2 => n17650, ZN => DataMem_N1663);
   U11692 : NOR2_X1 port map( A1 => n17006, A2 => n17661, ZN => DataMem_N2107);
   U11898 : NOR2_X1 port map( A1 => n17004, A2 => n17651, ZN => DataMem_N1727);
   U11726 : NOR2_X1 port map( A1 => n17006, A2 => n17658, ZN => DataMem_N2043);
   U11761 : NOR2_X1 port map( A1 => n17006, A2 => n17657, ZN => DataMem_N1979);
   U11863 : NOR2_X1 port map( A1 => n17004, A2 => n17654, ZN => DataMem_N1791);
   U11796 : NOR2_X1 port map( A1 => n17006, A2 => n17656, ZN => DataMem_N1915);
   U11830 : NOR2_X1 port map( A1 => n17006, A2 => n17655, ZN => DataMem_N1851);
   U11828 : NOR2_X1 port map( A1 => n17004, A2 => n17655, ZN => DataMem_N1855);
   U11865 : NOR2_X1 port map( A1 => n17006, A2 => n17654, ZN => DataMem_N1787);
   U11900 : NOR2_X1 port map( A1 => n17006, A2 => n17651, ZN => DataMem_N1723);
   U11794 : NOR2_X1 port map( A1 => n17004, A2 => n17656, ZN => DataMem_N1919);
   U11961 : NOR2_X1 port map( A1 => n17006, A2 => n17650, ZN => DataMem_N1659);
   U11635 : AOI22_X1 port map( A1 => n16823, A2 => DataMem_Mem_7_5_port, B1 => 
                           n17530, B2 => DataMem_Mem_6_5_port, ZN => n16951);
   U11634 : AOI22_X1 port map( A1 => n17531, A2 => DataMem_Mem_5_5_port, B1 => 
                           n16822, B2 => DataMem_Mem_4_5_port, ZN => n16952);
   U11633 : AOI22_X1 port map( A1 => n17122, A2 => DataMem_Mem_3_5_port, B1 => 
                           n17652, B2 => DataMem_Mem_2_5_port, ZN => n16953);
   U11632 : AOI22_X1 port map( A1 => n17124, A2 => DataMem_Mem_1_5_port, B1 => 
                           n16818, B2 => DataMem_Mem_0_5_port, ZN => n16954);
   U11630 : NOR2_X1 port map( A1 => n17155, A2 => n16950, ZN => DataMem_N2176);
   U11824 : NOR2_X1 port map( A1 => n17000, A2 => n16594, ZN => DataMem_N1863);
   U11790 : NOR2_X1 port map( A1 => n17000, A2 => n16593, ZN => DataMem_N1927);
   U11755 : NOR2_X1 port map( A1 => n17000, A2 => n16592, ZN => DataMem_N1991);
   U11720 : NOR2_X1 port map( A1 => n17000, A2 => n16591, ZN => DataMem_N2055);
   U11686 : NOR2_X1 port map( A1 => n17000, A2 => n16590, ZN => DataMem_N2119);
   U11611 : AOI22_X1 port map( A1 => n17660, A2 => DataMem_Mem_7_9_port, B1 => 
                           n16824, B2 => DataMem_Mem_6_9_port, ZN => n16931);
   U11610 : AOI22_X1 port map( A1 => n16821, A2 => DataMem_Mem_5_9_port, B1 => 
                           n16822, B2 => DataMem_Mem_4_9_port, ZN => n16932);
   U11609 : AOI22_X1 port map( A1 => n17122, A2 => DataMem_Mem_3_9_port, B1 => 
                           n17653, B2 => DataMem_Mem_2_9_port, ZN => n16933);
   U11608 : AOI22_X1 port map( A1 => n17124, A2 => DataMem_Mem_1_9_port, B1 => 
                           n16818, B2 => DataMem_Mem_0_9_port, ZN => n16934);
   U11606 : NOR2_X1 port map( A1 => n17155, A2 => n16930, ZN => DataMem_N2188);
   U11953 : NOR2_X1 port map( A1 => n17002, A2 => n16597, ZN => DataMem_N1667);
   U11896 : NOR2_X1 port map( A1 => n17002, A2 => n16596, ZN => DataMem_N1731);
   U11861 : NOR2_X1 port map( A1 => n17002, A2 => n16595, ZN => DataMem_N1795);
   U11826 : NOR2_X1 port map( A1 => n17002, A2 => n16594, ZN => DataMem_N1859);
   U11792 : NOR2_X1 port map( A1 => n17002, A2 => n16593, ZN => DataMem_N1923);
   U11757 : NOR2_X1 port map( A1 => n17002, A2 => n16592, ZN => DataMem_N1987);
   U11722 : NOR2_X1 port map( A1 => n17002, A2 => n16591, ZN => DataMem_N2051);
   U11688 : NOR2_X1 port map( A1 => n17002, A2 => n16590, ZN => DataMem_N2115);
   U11969 : NOR2_X1 port map( A1 => n17010, A2 => n17650, ZN => DataMem_N1651);
   U11659 : AOI22_X1 port map( A1 => n17659, A2 => DataMem_Mem_7_1_port, B1 => 
                           n17530, B2 => DataMem_Mem_6_1_port, ZN => n16971);
   U11658 : AOI22_X1 port map( A1 => n17531, A2 => DataMem_Mem_5_1_port, B1 => 
                           n16822, B2 => DataMem_Mem_4_1_port, ZN => n16972);
   U11657 : AOI22_X1 port map( A1 => n17122, A2 => DataMem_Mem_3_1_port, B1 => 
                           n17653, B2 => DataMem_Mem_2_1_port, ZN => n16973);
   U11656 : AOI22_X1 port map( A1 => n17124, A2 => DataMem_Mem_1_1_port, B1 => 
                           n17125, B2 => DataMem_Mem_0_1_port, ZN => n16974);
   U11654 : NOR2_X1 port map( A1 => n17155, A2 => n16970, ZN => DataMem_N2164);
   U11959 : NOR2_X1 port map( A1 => n17005, A2 => n17650, ZN => DataMem_N1661);
   U11629 : AOI22_X1 port map( A1 => n16823, A2 => DataMem_Mem_7_6_port, B1 => 
                           n17530, B2 => DataMem_Mem_6_6_port, ZN => n16946);
   U11628 : AOI22_X1 port map( A1 => n17531, A2 => DataMem_Mem_5_6_port, B1 => 
                           n16822, B2 => DataMem_Mem_4_6_port, ZN => n16947);
   U11627 : AOI22_X1 port map( A1 => n16819, A2 => DataMem_Mem_3_6_port, B1 => 
                           n17652, B2 => DataMem_Mem_2_6_port, ZN => n16948);
   U11626 : AOI22_X1 port map( A1 => n17124, A2 => DataMem_Mem_1_6_port, B1 => 
                           n17125, B2 => DataMem_Mem_0_6_port, ZN => n16949);
   U11624 : NOR2_X1 port map( A1 => n17155, A2 => n16945, ZN => DataMem_N2179);
   U11690 : NOR2_X1 port map( A1 => n17004, A2 => n17661, ZN => DataMem_N2111);
   U11771 : NOR2_X1 port map( A1 => n16981, A2 => n17656, ZN => DataMem_N1965);
   U11897 : NOR2_X1 port map( A1 => n17003, A2 => n16596, ZN => DataMem_N1729);
   U11736 : NOR2_X1 port map( A1 => n16981, A2 => n17657, ZN => DataMem_N2029);
   U11701 : NOR2_X1 port map( A1 => n16981, A2 => n17658, ZN => DataMem_N2093);
   U11667 : NOR2_X1 port map( A1 => n16981, A2 => n17661, ZN => DataMem_N2157);
   U11955 : NOR2_X1 port map( A1 => n17003, A2 => n16597, ZN => DataMem_N1665);
   U11491 : AOI22_X1 port map( A1 => n16823, A2 => DataMem_Mem_7_29_port, B1 =>
                           n16824, B2 => DataMem_Mem_6_29_port, ZN => n16831);
   U11490 : AOI22_X1 port map( A1 => n17531, A2 => DataMem_Mem_5_29_port, B1 =>
                           n16822, B2 => DataMem_Mem_4_29_port, ZN => n16832);
   U11489 : AOI22_X1 port map( A1 => n17122, A2 => DataMem_Mem_3_29_port, B1 =>
                           n17653, B2 => DataMem_Mem_2_29_port, ZN => n16833);
   U11488 : AOI22_X1 port map( A1 => n16817, A2 => DataMem_Mem_1_29_port, B1 =>
                           n17125, B2 => DataMem_Mem_0_29_port, ZN => n16834);
   U11486 : NOR2_X1 port map( A1 => n17155, A2 => n16830, ZN => DataMem_N2248);
   U11913 : NOR2_X1 port map( A1 => n16982, A2 => n17650, ZN => DataMem_N1707);
   U11617 : AOI22_X1 port map( A1 => n17659, A2 => DataMem_Mem_7_8_port, B1 => 
                           n16824, B2 => DataMem_Mem_6_8_port, ZN => n16936);
   U11616 : AOI22_X1 port map( A1 => n17531, A2 => DataMem_Mem_5_8_port, B1 => 
                           n16822, B2 => DataMem_Mem_4_8_port, ZN => n16937);
   U11615 : AOI22_X1 port map( A1 => n17122, A2 => DataMem_Mem_3_8_port, B1 => 
                           n17653, B2 => DataMem_Mem_2_8_port, ZN => n16938);
   U11614 : AOI22_X1 port map( A1 => n16817, A2 => DataMem_Mem_1_8_port, B1 => 
                           n16818, B2 => DataMem_Mem_0_8_port, ZN => n16939);
   U11612 : NOR2_X1 port map( A1 => n17155, A2 => n16935, ZN => DataMem_N2185);
   U11876 : NOR2_X1 port map( A1 => n16982, A2 => n17651, ZN => DataMem_N1771);
   U11841 : NOR2_X1 port map( A1 => n16982, A2 => n17654, ZN => DataMem_N1835);
   U11806 : NOR2_X1 port map( A1 => n16982, A2 => n17655, ZN => DataMem_N1899);
   U11772 : NOR2_X1 port map( A1 => n16982, A2 => n17656, ZN => DataMem_N1963);
   U11697 : NOR2_X1 port map( A1 => n17011, A2 => n17661, ZN => DataMem_N2097);
   U11737 : NOR2_X1 port map( A1 => n16982, A2 => n17657, ZN => DataMem_N2027);
   U11702 : NOR2_X1 port map( A1 => n16982, A2 => n17658, ZN => DataMem_N2091);
   U11668 : NOR2_X1 port map( A1 => n16982, A2 => n17661, ZN => DataMem_N2155);
   U11731 : NOR2_X1 port map( A1 => n17011, A2 => n17658, ZN => DataMem_N2033);
   U11503 : AOI22_X1 port map( A1 => n16823, A2 => DataMem_Mem_7_27_port, B1 =>
                           n17530, B2 => DataMem_Mem_6_27_port, ZN => n16841);
   U11502 : AOI22_X1 port map( A1 => n17531, A2 => DataMem_Mem_5_27_port, B1 =>
                           n16822, B2 => DataMem_Mem_4_27_port, ZN => n16842);
   U11501 : AOI22_X1 port map( A1 => n17122, A2 => DataMem_Mem_3_27_port, B1 =>
                           n17653, B2 => DataMem_Mem_2_27_port, ZN => n16843);
   U11500 : AOI22_X1 port map( A1 => n17124, A2 => DataMem_Mem_1_27_port, B1 =>
                           n17125, B2 => DataMem_Mem_0_27_port, ZN => n16844);
   U11498 : NOR2_X1 port map( A1 => n17155, A2 => n16840, ZN => DataMem_N2242);
   U11918 : AOI22_X1 port map( A1 => pipeline_Forward_sw1_mux, A2 => 
                           pipeline_data_to_RF_from_WB_27_port, B1 => n13793, 
                           B2 => n17743, ZN => n16984);
   U11917 : NOR2_X1 port map( A1 => n16984, A2 => n17650, ZN => DataMem_N1703);
   U11878 : NOR2_X1 port map( A1 => n16984, A2 => n17651, ZN => DataMem_N1767);
   U11766 : NOR2_X1 port map( A1 => n17011, A2 => n17657, ZN => DataMem_N1969);
   U11843 : NOR2_X1 port map( A1 => n16984, A2 => n17654, ZN => DataMem_N1831);
   U11808 : NOR2_X1 port map( A1 => n16984, A2 => n17655, ZN => DataMem_N1895);
   U11774 : NOR2_X1 port map( A1 => n16984, A2 => n17656, ZN => DataMem_N1959);
   U11801 : NOR2_X1 port map( A1 => n17011, A2 => n17656, ZN => DataMem_N1905);
   U11739 : NOR2_X1 port map( A1 => n16984, A2 => n17657, ZN => DataMem_N2023);
   U11672 : NOR2_X1 port map( A1 => n16986, A2 => n16590, ZN => DataMem_N2147);
   U11704 : NOR2_X1 port map( A1 => n16984, A2 => n17658, ZN => DataMem_N2087);
   U11670 : NOR2_X1 port map( A1 => n16984, A2 => n17661, ZN => DataMem_N2151);
   U11835 : NOR2_X1 port map( A1 => n17011, A2 => n17655, ZN => DataMem_N1841);
   U11509 : AOI22_X1 port map( A1 => n17660, A2 => DataMem_Mem_7_26_port, B1 =>
                           n17530, B2 => DataMem_Mem_6_26_port, ZN => n16846);
   U11508 : AOI22_X1 port map( A1 => n17531, A2 => DataMem_Mem_5_26_port, B1 =>
                           n16822, B2 => DataMem_Mem_4_26_port, ZN => n16847);
   U11507 : AOI22_X1 port map( A1 => n17122, A2 => DataMem_Mem_3_26_port, B1 =>
                           n17652, B2 => DataMem_Mem_2_26_port, ZN => n16848);
   U11506 : AOI22_X1 port map( A1 => n17124, A2 => DataMem_Mem_1_26_port, B1 =>
                           n17125, B2 => DataMem_Mem_0_26_port, ZN => n16849);
   U11504 : NOR2_X1 port map( A1 => n17155, A2 => n16845, ZN => DataMem_N2239);
   U11920 : AOI22_X1 port map( A1 => pipeline_Forward_sw1_mux, A2 => 
                           pipeline_data_to_RF_from_WB_26_port, B1 => n13794, 
                           B2 => n17380, ZN => n16985);
   U11919 : NOR2_X1 port map( A1 => n16985, A2 => n17650, ZN => DataMem_N1701);
   U11870 : NOR2_X1 port map( A1 => n17011, A2 => n17654, ZN => DataMem_N1777);
   U11879 : NOR2_X1 port map( A1 => n16985, A2 => n17651, ZN => DataMem_N1765);
   U11844 : NOR2_X1 port map( A1 => n16985, A2 => n17654, ZN => DataMem_N1829);
   U11809 : NOR2_X1 port map( A1 => n16985, A2 => n17655, ZN => DataMem_N1893);
   U11905 : NOR2_X1 port map( A1 => n17011, A2 => n17651, ZN => DataMem_N1713);
   U11775 : NOR2_X1 port map( A1 => n16985, A2 => n17656, ZN => DataMem_N1957);
   U11740 : NOR2_X1 port map( A1 => n16985, A2 => n17657, ZN => DataMem_N2021);
   U11705 : NOR2_X1 port map( A1 => n16985, A2 => n17658, ZN => DataMem_N2085);
   U11971 : NOR2_X1 port map( A1 => n17011, A2 => n17650, ZN => DataMem_N1649);
   U11671 : NOR2_X1 port map( A1 => n16985, A2 => n17661, ZN => DataMem_N2149);
   U11665 : AOI22_X1 port map( A1 => n17659, A2 => DataMem_Mem_7_0_port, B1 => 
                           n17530, B2 => DataMem_Mem_6_0_port, ZN => n16976);
   U11664 : AOI22_X1 port map( A1 => n17531, A2 => DataMem_Mem_5_0_port, B1 => 
                           n16822, B2 => DataMem_Mem_4_0_port, ZN => n16977);
   U11663 : AOI22_X1 port map( A1 => n17122, A2 => DataMem_Mem_3_0_port, B1 => 
                           n17652, B2 => DataMem_Mem_2_0_port, ZN => n16978);
   U11662 : AOI22_X1 port map( A1 => n17124, A2 => DataMem_Mem_1_0_port, B1 => 
                           n17125, B2 => DataMem_Mem_0_0_port, ZN => n16979);
   U11660 : NOR2_X1 port map( A1 => n17155, A2 => n16975, ZN => DataMem_N2161);
   U11515 : AOI22_X1 port map( A1 => n17660, A2 => DataMem_Mem_7_25_port, B1 =>
                           n17530, B2 => DataMem_Mem_6_25_port, ZN => n16851);
   U11514 : AOI22_X1 port map( A1 => n17531, A2 => DataMem_Mem_5_25_port, B1 =>
                           n16822, B2 => DataMem_Mem_4_25_port, ZN => n16852);
   U11513 : AOI22_X1 port map( A1 => n17122, A2 => DataMem_Mem_3_25_port, B1 =>
                           n16820, B2 => DataMem_Mem_2_25_port, ZN => n16853);
   U11512 : AOI22_X1 port map( A1 => n17124, A2 => DataMem_Mem_1_25_port, B1 =>
                           n16818, B2 => DataMem_Mem_0_25_port, ZN => n16854);
   U11510 : NOR2_X1 port map( A1 => n17155, A2 => n16850, ZN => DataMem_N2236);
   U11921 : NOR2_X1 port map( A1 => n16986, A2 => n16597, ZN => DataMem_N1699);
   U11880 : NOR2_X1 port map( A1 => n16986, A2 => n16596, ZN => DataMem_N1763);
   U11910 : AOI22_X1 port map( A1 => pipeline_Forward_sw1_mux, A2 => 
                           pipeline_data_to_RF_from_WB_31_port, B1 => n13783, 
                           B2 => n17380, ZN => n16980);
   U11700 : NOR2_X1 port map( A1 => n16980, A2 => n17658, ZN => DataMem_N2095);
   U11845 : NOR2_X1 port map( A1 => n16986, A2 => n16595, ZN => DataMem_N1827);
   U11810 : NOR2_X1 port map( A1 => n16986, A2 => n16594, ZN => DataMem_N1891);
   U11735 : NOR2_X1 port map( A1 => n16980, A2 => n17657, ZN => DataMem_N2031);
   U11776 : NOR2_X1 port map( A1 => n16986, A2 => n16593, ZN => DataMem_N1955);
   U11741 : NOR2_X1 port map( A1 => n16986, A2 => n16592, ZN => DataMem_N2019);
   U11706 : NOR2_X1 port map( A1 => n16986, A2 => n16591, ZN => DataMem_N2083);
   U11770 : NOR2_X1 port map( A1 => n16980, A2 => n17656, ZN => DataMem_N1967);
   U11915 : NOR2_X1 port map( A1 => n16983, A2 => n17650, ZN => DataMem_N1705);
   U11877 : NOR2_X1 port map( A1 => n16983, A2 => n17651, ZN => DataMem_N1769);
   U11673 : NOR2_X1 port map( A1 => n16987, A2 => n16590, ZN => DataMem_N2145);
   U11842 : NOR2_X1 port map( A1 => n16983, A2 => n17654, ZN => DataMem_N1833);
   U11807 : NOR2_X1 port map( A1 => n16983, A2 => n17655, ZN => DataMem_N1897);
   U11773 : NOR2_X1 port map( A1 => n16983, A2 => n17656, ZN => DataMem_N1961);
   U11707 : NOR2_X1 port map( A1 => n16987, A2 => n16591, ZN => DataMem_N2081);
   U11738 : NOR2_X1 port map( A1 => n16983, A2 => n17657, ZN => DataMem_N2025);
   U11703 : NOR2_X1 port map( A1 => n16983, A2 => n17658, ZN => DataMem_N2089);
   U11742 : NOR2_X1 port map( A1 => n16987, A2 => n16592, ZN => DataMem_N2017);
   U11669 : NOR2_X1 port map( A1 => n16983, A2 => n17661, ZN => DataMem_N2153);
   U11581 : AOI22_X1 port map( A1 => n17659, A2 => DataMem_Mem_7_14_port, B1 =>
                           n17530, B2 => DataMem_Mem_6_14_port, ZN => n16906);
   U11580 : AOI22_X1 port map( A1 => n16821, A2 => DataMem_Mem_5_14_port, B1 =>
                           n16822, B2 => DataMem_Mem_4_14_port, ZN => n16907);
   U11579 : AOI22_X1 port map( A1 => n17122, A2 => DataMem_Mem_3_14_port, B1 =>
                           n17653, B2 => DataMem_Mem_2_14_port, ZN => n16908);
   U11578 : AOI22_X1 port map( A1 => n17124, A2 => DataMem_Mem_1_14_port, B1 =>
                           n16818, B2 => DataMem_Mem_0_14_port, ZN => n16909);
   U11576 : NOR2_X1 port map( A1 => n17155, A2 => n16905, ZN => DataMem_N2203);
   U11943 : NOR2_X1 port map( A1 => n16997, A2 => n17650, ZN => DataMem_N1677);
   U11891 : NOR2_X1 port map( A1 => n16997, A2 => n17651, ZN => DataMem_N1741);
   U11777 : NOR2_X1 port map( A1 => n16987, A2 => n16593, ZN => DataMem_N1953);
   U11856 : NOR2_X1 port map( A1 => n16997, A2 => n17654, ZN => DataMem_N1805);
   U11821 : NOR2_X1 port map( A1 => n16997, A2 => n17655, ZN => DataMem_N1869);
   U11787 : NOR2_X1 port map( A1 => n16997, A2 => n17656, ZN => DataMem_N1933);
   U11811 : NOR2_X1 port map( A1 => n16987, A2 => n16594, ZN => DataMem_N1889);
   U11752 : NOR2_X1 port map( A1 => n16997, A2 => n17657, ZN => DataMem_N1997);
   U11717 : NOR2_X1 port map( A1 => n16997, A2 => n17658, ZN => DataMem_N2061);
   U11846 : NOR2_X1 port map( A1 => n16987, A2 => n16595, ZN => DataMem_N1825);
   U11683 : NOR2_X1 port map( A1 => n16997, A2 => n17661, ZN => DataMem_N2125);
   U11575 : AOI22_X1 port map( A1 => n17659, A2 => DataMem_Mem_7_15_port, B1 =>
                           n16824, B2 => DataMem_Mem_6_15_port, ZN => n16901);
   U11574 : AOI22_X1 port map( A1 => n16821, A2 => DataMem_Mem_5_15_port, B1 =>
                           n16822, B2 => DataMem_Mem_4_15_port, ZN => n16902);
   U11573 : AOI22_X1 port map( A1 => n17122, A2 => DataMem_Mem_3_15_port, B1 =>
                           n17653, B2 => DataMem_Mem_2_15_port, ZN => n16903);
   U11572 : AOI22_X1 port map( A1 => n16817, A2 => DataMem_Mem_1_15_port, B1 =>
                           n17125, B2 => DataMem_Mem_0_15_port, ZN => n16904);
   U11570 : NOR2_X1 port map( A1 => n12766, A2 => n16900, ZN => DataMem_N2206);
   U11881 : NOR2_X1 port map( A1 => n16987, A2 => n16596, ZN => DataMem_N1761);
   U11941 : NOR2_X1 port map( A1 => n16996, A2 => n17650, ZN => DataMem_N1679);
   U11890 : NOR2_X1 port map( A1 => n16996, A2 => n17651, ZN => DataMem_N1743);
   U11855 : NOR2_X1 port map( A1 => n16996, A2 => n17654, ZN => DataMem_N1807);
   U11923 : NOR2_X1 port map( A1 => n16987, A2 => n16597, ZN => DataMem_N1697);
   U11820 : NOR2_X1 port map( A1 => n16996, A2 => n17655, ZN => DataMem_N1871);
   U11521 : AOI22_X1 port map( A1 => n17660, A2 => DataMem_Mem_7_24_port, B1 =>
                           n17530, B2 => DataMem_Mem_6_24_port, ZN => n16856);
   U11520 : AOI22_X1 port map( A1 => n17531, A2 => DataMem_Mem_5_24_port, B1 =>
                           n16822, B2 => DataMem_Mem_4_24_port, ZN => n16857);
   U11519 : AOI22_X1 port map( A1 => n16819, A2 => DataMem_Mem_3_24_port, B1 =>
                           n16820, B2 => DataMem_Mem_2_24_port, ZN => n16858);
   U11518 : AOI22_X1 port map( A1 => n16817, A2 => DataMem_Mem_1_24_port, B1 =>
                           n16818, B2 => DataMem_Mem_0_24_port, ZN => n16859);
   U11516 : NOR2_X1 port map( A1 => n17155, A2 => n16855, ZN => DataMem_N2233);
   U11786 : NOR2_X1 port map( A1 => n16996, A2 => n17656, ZN => DataMem_N1935);
   U11751 : NOR2_X1 port map( A1 => n16996, A2 => n17657, ZN => DataMem_N1999);
   U11716 : NOR2_X1 port map( A1 => n16996, A2 => n17658, ZN => DataMem_N2063);
   U11689 : NOR2_X1 port map( A1 => n17003, A2 => n16590, ZN => DataMem_N2113);
   U11682 : NOR2_X1 port map( A1 => n16996, A2 => n17661, ZN => DataMem_N2127);
   U11587 : AOI22_X1 port map( A1 => n17659, A2 => DataMem_Mem_7_13_port, B1 =>
                           n16824, B2 => DataMem_Mem_6_13_port, ZN => n16911);
   U11586 : AOI22_X1 port map( A1 => n16821, A2 => DataMem_Mem_5_13_port, B1 =>
                           n16822, B2 => DataMem_Mem_4_13_port, ZN => n16912);
   U11585 : AOI22_X1 port map( A1 => n17122, A2 => DataMem_Mem_3_13_port, B1 =>
                           n17653, B2 => DataMem_Mem_2_13_port, ZN => n16913);
   U11584 : AOI22_X1 port map( A1 => n16817, A2 => DataMem_Mem_1_13_port, B1 =>
                           n17125, B2 => DataMem_Mem_0_13_port, ZN => n16914);
   U11582 : NOR2_X1 port map( A1 => n12766, A2 => n16910, ZN => DataMem_N2200);
   U11946 : AOI22_X1 port map( A1 => pipeline_Forward_sw1_mux, A2 => 
                           pipeline_data_to_RF_from_WB_13_port, B1 => n13790, 
                           B2 => n17380, ZN => n16998);
   U11945 : NOR2_X1 port map( A1 => n16998, A2 => n17650, ZN => DataMem_N1675);
   U11723 : NOR2_X1 port map( A1 => n17003, A2 => n16591, ZN => DataMem_N2049);
   U11892 : NOR2_X1 port map( A1 => n16998, A2 => n17651, ZN => DataMem_N1739);
   U11857 : NOR2_X1 port map( A1 => n16998, A2 => n17654, ZN => DataMem_N1803);
   U11758 : NOR2_X1 port map( A1 => n17003, A2 => n16592, ZN => DataMem_N1985);
   U11822 : NOR2_X1 port map( A1 => n16998, A2 => n17655, ZN => DataMem_N1867);
   U11788 : NOR2_X1 port map( A1 => n16998, A2 => n17656, ZN => DataMem_N1931);
   U11753 : NOR2_X1 port map( A1 => n16998, A2 => n17657, ZN => DataMem_N1995);
   U11793 : NOR2_X1 port map( A1 => n17003, A2 => n16593, ZN => DataMem_N1921);
   U11718 : NOR2_X1 port map( A1 => n16998, A2 => n17658, ZN => DataMem_N2059);
   U11684 : NOR2_X1 port map( A1 => n16998, A2 => n17661, ZN => DataMem_N2123);
   U11827 : NOR2_X1 port map( A1 => n17003, A2 => n16594, ZN => DataMem_N1857);
   U11485 : AOI22_X1 port map( A1 => n17659, A2 => DataMem_Mem_7_30_port, B1 =>
                           n16824, B2 => DataMem_Mem_6_30_port, ZN => n16826);
   U11484 : AOI22_X1 port map( A1 => n17531, A2 => DataMem_Mem_5_30_port, B1 =>
                           n16822, B2 => DataMem_Mem_4_30_port, ZN => n16827);
   U11483 : AOI22_X1 port map( A1 => n17122, A2 => DataMem_Mem_3_30_port, B1 =>
                           n17653, B2 => DataMem_Mem_2_30_port, ZN => n16828);
   U11482 : AOI22_X1 port map( A1 => n17124, A2 => DataMem_Mem_1_30_port, B1 =>
                           n16818, B2 => DataMem_Mem_0_30_port, ZN => n16829);
   U11480 : NOR2_X1 port map( A1 => n17155, A2 => n16825, ZN => DataMem_N2251);
   U11911 : NOR2_X1 port map( A1 => n16981, A2 => n17650, ZN => DataMem_N1709);
   U11875 : NOR2_X1 port map( A1 => n16981, A2 => n17651, ZN => DataMem_N1773);
   U11840 : NOR2_X1 port map( A1 => n16981, A2 => n17654, ZN => DataMem_N1837);
   U11862 : NOR2_X1 port map( A1 => n17003, A2 => n16595, ZN => DataMem_N1793);
   U11805 : NOR2_X1 port map( A1 => n16981, A2 => n17655, ZN => DataMem_N1901);
   U11724 : NOR2_X1 port map( A1 => n17004, A2 => n17658, ZN => DataMem_N2047);
   U11497 : AOI22_X1 port map( A1 => n16823, A2 => DataMem_Mem_7_28_port, B1 =>
                           n17530, B2 => DataMem_Mem_6_28_port, ZN => n16836);
   U11496 : AOI22_X1 port map( A1 => n17531, A2 => DataMem_Mem_5_28_port, B1 =>
                           n16822, B2 => DataMem_Mem_4_28_port, ZN => n16837);
   U11495 : AOI22_X1 port map( A1 => n17122, A2 => DataMem_Mem_3_28_port, B1 =>
                           n17653, B2 => DataMem_Mem_2_28_port, ZN => n16838);
   U11494 : AOI22_X1 port map( A1 => n17124, A2 => DataMem_Mem_1_28_port, B1 =>
                           n17125, B2 => DataMem_Mem_0_28_port, ZN => n16839);
   U11492 : NOR2_X1 port map( A1 => n12766, A2 => n16835, ZN => DataMem_N2245);
   U11710 : NOR2_X1 port map( A1 => n16990, A2 => n16591, ZN => DataMem_N2075);
   U11818 : NOR2_X1 port map( A1 => n16994, A2 => n16594, ZN => DataMem_N1875);
   U11676 : NOR2_X1 port map( A1 => n16990, A2 => n16590, ZN => DataMem_N2139);
   U11545 : AOI22_X1 port map( A1 => n17660, A2 => DataMem_Mem_7_20_port, B1 =>
                           n17530, B2 => DataMem_Mem_6_20_port, ZN => n16876);
   U11544 : AOI22_X1 port map( A1 => n16821, A2 => DataMem_Mem_5_20_port, B1 =>
                           n16822, B2 => DataMem_Mem_4_20_port, ZN => n16877);
   U11543 : AOI22_X1 port map( A1 => n16819, A2 => DataMem_Mem_3_20_port, B1 =>
                           n17653, B2 => DataMem_Mem_2_20_port, ZN => n16878);
   U11542 : AOI22_X1 port map( A1 => n17124, A2 => DataMem_Mem_1_20_port, B1 =>
                           n17125, B2 => DataMem_Mem_0_20_port, ZN => n16879);
   U11540 : NOR2_X1 port map( A1 => n17155, A2 => n16875, ZN => DataMem_N2221);
   U11931 : NOR2_X1 port map( A1 => n16991, A2 => n16597, ZN => DataMem_N1689);
   U11885 : NOR2_X1 port map( A1 => n16991, A2 => n16596, ZN => DataMem_N1753);
   U11850 : NOR2_X1 port map( A1 => n16991, A2 => n16595, ZN => DataMem_N1817);
   U11815 : NOR2_X1 port map( A1 => n16991, A2 => n16594, ZN => DataMem_N1881);
   U11781 : NOR2_X1 port map( A1 => n16991, A2 => n16593, ZN => DataMem_N1945);
   U11853 : NOR2_X1 port map( A1 => n16994, A2 => n16595, ZN => DataMem_N1811);
   U11746 : NOR2_X1 port map( A1 => n16991, A2 => n16592, ZN => DataMem_N2009);
   U11711 : NOR2_X1 port map( A1 => n16991, A2 => n16591, ZN => DataMem_N2073);
   U11677 : NOR2_X1 port map( A1 => n16991, A2 => n16590, ZN => DataMem_N2137);
   U11551 : AOI22_X1 port map( A1 => n17659, A2 => DataMem_Mem_7_19_port, B1 =>
                           n16824, B2 => DataMem_Mem_6_19_port, ZN => n16881);
   U11550 : AOI22_X1 port map( A1 => n16821, A2 => DataMem_Mem_5_19_port, B1 =>
                           n16822, B2 => DataMem_Mem_4_19_port, ZN => n16882);
   U11549 : AOI22_X1 port map( A1 => n17122, A2 => DataMem_Mem_3_19_port, B1 =>
                           n16820, B2 => DataMem_Mem_2_19_port, ZN => n16883);
   U11548 : AOI22_X1 port map( A1 => n17124, A2 => DataMem_Mem_1_19_port, B1 =>
                           n16818, B2 => DataMem_Mem_0_19_port, ZN => n16884);
   U11546 : NOR2_X1 port map( A1 => n17155, A2 => n16880, ZN => DataMem_N2218);
   U11888 : NOR2_X1 port map( A1 => n16994, A2 => n16596, ZN => DataMem_N1747);
   U11934 : AOI22_X1 port map( A1 => pipeline_Forward_sw1_mux, A2 => 
                           pipeline_data_to_RF_from_WB_19_port, B1 => n13800, 
                           B2 => n17380, ZN => n16992);
   U11933 : NOR2_X1 port map( A1 => n16992, A2 => n16597, ZN => DataMem_N1687);
   U11886 : NOR2_X1 port map( A1 => n16992, A2 => n16596, ZN => DataMem_N1751);
   U11936 : AOI22_X1 port map( A1 => pipeline_Forward_sw1_mux, A2 => 
                           pipeline_data_to_RF_from_WB_18_port, B1 => n13801, 
                           B2 => n17380, ZN => n16993);
   U11713 : NOR2_X1 port map( A1 => n16993, A2 => n16591, ZN => DataMem_N2069);
   U11851 : NOR2_X1 port map( A1 => n16992, A2 => n16595, ZN => DataMem_N1815);
   U11816 : NOR2_X1 port map( A1 => n16992, A2 => n16594, ZN => DataMem_N1879);
   U11937 : NOR2_X1 port map( A1 => n16994, A2 => n16597, ZN => DataMem_N1683);
   U11782 : NOR2_X1 port map( A1 => n16992, A2 => n16593, ZN => DataMem_N1943);
   U11563 : AOI22_X1 port map( A1 => n17660, A2 => DataMem_Mem_7_17_port, B1 =>
                           n16824, B2 => DataMem_Mem_6_17_port, ZN => n16891);
   U11562 : AOI22_X1 port map( A1 => n16821, A2 => DataMem_Mem_5_17_port, B1 =>
                           n16822, B2 => DataMem_Mem_4_17_port, ZN => n16892);
   U11561 : AOI22_X1 port map( A1 => n17122, A2 => DataMem_Mem_3_17_port, B1 =>
                           n16820, B2 => DataMem_Mem_2_17_port, ZN => n16893);
   U11560 : AOI22_X1 port map( A1 => n17124, A2 => DataMem_Mem_1_17_port, B1 =>
                           n17125, B2 => DataMem_Mem_0_17_port, ZN => n16894);
   U11558 : NOR2_X1 port map( A1 => n17155, A2 => n16890, ZN => DataMem_N2212);
   U11747 : NOR2_X1 port map( A1 => n16992, A2 => n16592, ZN => DataMem_N2007);
   U8521 : NAND4_X1 port map( A1 => n14116, A2 => n14117, A3 => n14113, A4 => 
                           n14100, ZN => n14121);
   U8520 : NOR2_X1 port map( A1 => n14120, A2 => n14121, ZN => n14096);
   U8508 : NOR4_X1 port map( A1 => n14096, A2 => n14097, A3 => n14098, A4 => 
                           n14099, ZN => n14095);
   U8519 : AOI22_X1 port map( A1 => 
                           pipeline_stageD_offset_jump_sign_ext_21_port, A2 => 
                           n14116, B1 => 
                           pipeline_stageD_offset_jump_sign_ext_22_port, B2 => 
                           n14117, ZN => n14119);
   U8518 : OAI221_X1 port map( B1 => 
                           pipeline_stageD_offset_jump_sign_ext_21_port, B2 => 
                           n14116, C1 => 
                           pipeline_stageD_offset_jump_sign_ext_22_port, C2 => 
                           n14117, A => n14119, ZN => n14087);
   U8526 : NAND2_X1 port map( A1 => n14123, A2 => n17704, ZN => n13983);
   U8527 : NOR2_X1 port map( A1 => n17449, A2 => n14122, ZN => n14093);
   U8507 : AOI22_X1 port map( A1 => n14091, A2 => n14092, B1 => n14093, B2 => 
                           n14094, ZN => n14088);
   U8524 : NOR2_X1 port map( A1 => n14091, A2 => n14122, ZN => n14090);
   U8506 : OAI211_X1 port map( C1 => n14086, C2 => n14087, A => n14088, B => 
                           n14089, ZN => pipeline_cu_hazard_N40);
   U11712 : NOR2_X1 port map( A1 => n16992, A2 => n16591, ZN => DataMem_N2071);
   U8467 : OAI21_X1 port map( B1 => n14031, B2 => n14032, A => n14033, ZN => 
                           n14013);
   U8491 : NAND2_X1 port map( A1 => n14005, A2 => n13990, ZN => n14030);
   U8465 : NOR3_X1 port map( A1 => n14027, A2 => n14015, A3 => n14007, ZN => 
                           n14026);
   U8464 : NAND4_X1 port map( A1 => n14025, A2 => n14013, A3 => n14002, A4 => 
                           n14026, ZN => pipeline_cu_pipeline_N105);
   U11678 : NOR2_X1 port map( A1 => n16992, A2 => n16590, ZN => DataMem_N2135);
   U8488 : NOR2_X1 port map( A1 => n17313, A2 => n14047, ZN => n14000);
   U8452 : OAI221_X1 port map( B1 => n13999, B2 => n14000, C1 => n13999, C2 => 
                           n14001, A => n17704, ZN => n13985);
   U8451 : NOR2_X1 port map( A1 => Rst, A2 => n13998, ZN => n13994);
   U8469 : NOR3_X1 port map( A1 => n17347, A2 => n17409, A3 => n17313, ZN => 
                           n13995);
   U8450 : OAI21_X1 port map( B1 => Rst, B2 => n13997, A => n13983, ZN => 
                           n13996);
   U8449 : AOI221_X1 port map( B1 => n13993, B2 => n13994, C1 => n13995, C2 => 
                           n13994, A => n13996, ZN => n13986);
   U8448 : NOR2_X1 port map( A1 => Rst, A2 => n13984, ZN => n13992);
   U8447 : OAI221_X1 port map( B1 => n13989, B2 => n13990, C1 => n13989, C2 => 
                           n17076, A => n13992, ZN => n13987);
   U8446 : NAND4_X1 port map( A1 => n13985, A2 => n13986, A3 => n13987, A4 => 
                           n13988, ZN => pipeline_cu_pipeline_N110);
   U11557 : AOI22_X1 port map( A1 => n17659, A2 => DataMem_Mem_7_18_port, B1 =>
                           n16824, B2 => DataMem_Mem_6_18_port, ZN => n16886);
   U11556 : AOI22_X1 port map( A1 => n16821, A2 => DataMem_Mem_5_18_port, B1 =>
                           n16822, B2 => DataMem_Mem_4_18_port, ZN => n16887);
   U11555 : AOI22_X1 port map( A1 => n16819, A2 => DataMem_Mem_3_18_port, B1 =>
                           n17653, B2 => DataMem_Mem_2_18_port, ZN => n16888);
   U11554 : AOI22_X1 port map( A1 => n16817, A2 => DataMem_Mem_1_18_port, B1 =>
                           n17125, B2 => DataMem_Mem_0_18_port, ZN => n16889);
   U11552 : NOR2_X1 port map( A1 => n12766, A2 => n16885, ZN => DataMem_N2215);
   U8442 : NAND2_X1 port map( A1 => n13980, A2 => n13981, ZN => 
                           pipeline_cu_pipeline_N88);
   U11935 : NOR2_X1 port map( A1 => n16993, A2 => n16597, ZN => DataMem_N1685);
   U8490 : NOR2_X1 port map( A1 => n14047, A2 => n14058, ZN => n14068);
   U8487 : OAI211_X1 port map( C1 => n14012, C2 => n14024, A => n14029, B => 
                           n14070, ZN => n14069);
   U8486 : NOR2_X1 port map( A1 => n14068, A2 => n14069, ZN => n14053);
   U8475 : OAI211_X1 port map( C1 => n17406, C2 => n14030, A => n14053, B => 
                           n14041, ZN => pipeline_cu_pipeline_N102);
   U11887 : NOR2_X1 port map( A1 => n16993, A2 => n16596, ZN => DataMem_N1749);
   U11679 : NOR2_X1 port map( A1 => n16993, A2 => n16590, ZN => DataMem_N2133);
   U8501 : OAI22_X1 port map( A1 => n13993, A2 => n17348, B1 => n14084, B2 => 
                           n17532, ZN => n14083);
   U8500 : AOI211_X1 port map( C1 => 
                           pipeline_stageD_offset_to_jump_temp_10_port, C2 => 
                           pipeline_cu_pipeline_N89, A => n14009, B => n14083, 
                           ZN => n14073);
   U8499 : AOI221_X1 port map( B1 => pipeline_inst_IFID_DEC_27_port, B2 => 
                           pipeline_inst_IFID_DEC_26_port, C1 => n17313, C2 => 
                           n13993, A => pipeline_inst_IFID_DEC_29_port, ZN => 
                           n14075);
   U8498 : OAI21_X1 port map( B1 => pipeline_stageD_offset_to_jump_temp_9_port,
                           B2 => pipeline_stageD_offset_to_jump_temp_8_port, A 
                           => pipeline_cu_pipeline_N89, ZN => n14082);
   U8497 : OAI211_X1 port map( C1 => pipeline_inst_IFID_DEC_29_port, C2 => 
                           n17348, A => n14082, B => n14058, ZN => n14076);
   U8495 : AOI21_X1 port map( B1 => n17361, B2 => n17412, A => n13984, ZN => 
                           n14077);
   U8494 : AOI21_X1 port map( B1 => pipeline_stageD_offset_to_jump_temp_5_port,
                           B2 => n17410, A => n13984, ZN => n14078);
   U8493 : NOR4_X1 port map( A1 => n14075, A2 => n14076, A3 => n14077, A4 => 
                           n14078, ZN => n14074);
   U8492 : NAND4_X1 port map( A1 => n14071, A2 => n14072, A3 => n14073, A4 => 
                           n14074, ZN => pipeline_cu_pipeline_N101);
   U11852 : NOR2_X1 port map( A1 => n16993, A2 => n16595, ZN => DataMem_N1813);
   U8463 : AOI21_X1 port map( B1 => n14023, B2 => n14024, A => n14012, ZN => 
                           n14010);
   U8461 : NAND4_X1 port map( A1 => n14018, A2 => n14019, A3 => n14020, A4 => 
                           n14021, ZN => n14017);
   U8460 : NOR4_X1 port map( A1 => n14015, A2 => n14016, A3 => n14010, A4 => 
                           n14017, ZN => n14014);
   U8459 : OAI211_X1 port map( C1 => n14006, C2 => n14012, A => n14013, B => 
                           n14014, ZN => pipeline_cu_pipeline_N106);
   U8468 : OAI211_X1 port map( C1 => n14023, C2 => n14012, A => n14034, B => 
                           n14035, ZN => pipeline_cu_pipeline_N104);
   U11817 : NOR2_X1 port map( A1 => n16993, A2 => n16594, ZN => DataMem_N1877);
   U8473 : OAI21_X1 port map( B1 => n14011, B2 => n14047, A => n14048, ZN => 
                           n14046);
   U8472 : AOI211_X1 port map( C1 => n14045, C2 => n14005, A => n14015, B => 
                           n14046, ZN => n14043);
   U8471 : NAND4_X1 port map( A1 => n14041, A2 => n14042, A3 => n14043, A4 => 
                           n14021, ZN => pipeline_cu_pipeline_N103);
   U11783 : NOR2_X1 port map( A1 => n16993, A2 => n16593, ZN => DataMem_N1941);
   U11748 : NOR2_X1 port map( A1 => n16993, A2 => n16592, ZN => DataMem_N2005);
   U11889 : NOR2_X1 port map( A1 => n16995, A2 => n17651, ZN => DataMem_N1745);
   U11527 : AOI22_X1 port map( A1 => n17660, A2 => DataMem_Mem_7_23_port, B1 =>
                           n17530, B2 => DataMem_Mem_6_23_port, ZN => n16861);
   U11526 : AOI22_X1 port map( A1 => n17531, A2 => DataMem_Mem_5_23_port, B1 =>
                           n16822, B2 => DataMem_Mem_4_23_port, ZN => n16862);
   U11525 : AOI22_X1 port map( A1 => n17122, A2 => DataMem_Mem_3_23_port, B1 =>
                           n16820, B2 => DataMem_Mem_2_23_port, ZN => n16863);
   U11524 : AOI22_X1 port map( A1 => n17124, A2 => DataMem_Mem_1_23_port, B1 =>
                           n17125, B2 => DataMem_Mem_0_23_port, ZN => n16864);
   U11522 : NOR2_X1 port map( A1 => n17155, A2 => n16860, ZN => DataMem_N2230);
   U11925 : NOR2_X1 port map( A1 => n16988, A2 => n16597, ZN => DataMem_N1695);
   U11804 : NOR2_X1 port map( A1 => n16980, A2 => n17655, ZN => DataMem_N1903);
   U11666 : NOR2_X1 port map( A1 => n16980, A2 => n17661, ZN => DataMem_N2159);
   U11882 : NOR2_X1 port map( A1 => n16988, A2 => n16596, ZN => DataMem_N1759);
   U11939 : NOR2_X1 port map( A1 => n16995, A2 => n17650, ZN => DataMem_N1681);
   U11847 : NOR2_X1 port map( A1 => n16988, A2 => n16595, ZN => DataMem_N1823);
   U11839 : NOR2_X1 port map( A1 => n16980, A2 => n17654, ZN => DataMem_N1839);
   U11479 : AOI22_X1 port map( A1 => n17659, A2 => DataMem_Mem_7_31_port, B1 =>
                           n16824, B2 => DataMem_Mem_6_31_port, ZN => n16813);
   U11478 : AOI22_X1 port map( A1 => n16821, A2 => DataMem_Mem_5_31_port, B1 =>
                           n16822, B2 => DataMem_Mem_4_31_port, ZN => n16814);
   U11477 : AOI22_X1 port map( A1 => n17122, A2 => DataMem_Mem_3_31_port, B1 =>
                           n17652, B2 => DataMem_Mem_2_31_port, ZN => n16815);
   U11476 : AOI22_X1 port map( A1 => n16817, A2 => DataMem_Mem_1_31_port, B1 =>
                           n17125, B2 => DataMem_Mem_0_31_port, ZN => n16816);
   U11474 : NOR2_X1 port map( A1 => n12766, A2 => n16812, ZN => DataMem_N2254);
   U11812 : NOR2_X1 port map( A1 => n16988, A2 => n16594, ZN => DataMem_N1887);
   U11569 : AOI22_X1 port map( A1 => n17659, A2 => DataMem_Mem_7_16_port, B1 =>
                           n16824, B2 => DataMem_Mem_6_16_port, ZN => n16896);
   U11568 : AOI22_X1 port map( A1 => n16821, A2 => DataMem_Mem_5_16_port, B1 =>
                           n16822, B2 => DataMem_Mem_4_16_port, ZN => n16897);
   U11567 : AOI22_X1 port map( A1 => n17122, A2 => DataMem_Mem_3_16_port, B1 =>
                           n17653, B2 => DataMem_Mem_2_16_port, ZN => n16898);
   U11566 : AOI22_X1 port map( A1 => n17124, A2 => DataMem_Mem_1_16_port, B1 =>
                           n17125, B2 => DataMem_Mem_0_16_port, ZN => n16899);
   U11564 : NOR2_X1 port map( A1 => n17155, A2 => n16895, ZN => DataMem_N2209);
   U11778 : NOR2_X1 port map( A1 => n16988, A2 => n16593, ZN => DataMem_N1951);
   U11874 : NOR2_X1 port map( A1 => n16980, A2 => n17651, ZN => DataMem_N1775);
   U11743 : NOR2_X1 port map( A1 => n16988, A2 => n16592, ZN => DataMem_N2015);
   U11708 : NOR2_X1 port map( A1 => n16988, A2 => n16591, ZN => DataMem_N2079);
   U11909 : NOR2_X1 port map( A1 => n16980, A2 => n17650, ZN => DataMem_N1711);
   U11674 : NOR2_X1 port map( A1 => n16988, A2 => n16590, ZN => DataMem_N2143);
   U11680 : NOR2_X1 port map( A1 => n16994, A2 => n16590, ZN => DataMem_N2131);
   U11533 : AOI22_X1 port map( A1 => n17660, A2 => DataMem_Mem_7_22_port, B1 =>
                           n17530, B2 => DataMem_Mem_6_22_port, ZN => n16866);
   U11532 : AOI22_X1 port map( A1 => n17531, A2 => DataMem_Mem_5_22_port, B1 =>
                           n16822, B2 => DataMem_Mem_4_22_port, ZN => n16867);
   U11531 : AOI22_X1 port map( A1 => n17122, A2 => DataMem_Mem_3_22_port, B1 =>
                           n16820, B2 => DataMem_Mem_2_22_port, ZN => n16868);
   U11530 : AOI22_X1 port map( A1 => n17124, A2 => DataMem_Mem_1_22_port, B1 =>
                           n17125, B2 => DataMem_Mem_0_22_port, ZN => n16869);
   U11528 : NOR2_X1 port map( A1 => n17155, A2 => n16865, ZN => DataMem_N2227);
   U11928 : AOI22_X1 port map( A1 => pipeline_Forward_sw1_mux, A2 => 
                           pipeline_data_to_RF_from_WB_22_port, B1 => n13797, 
                           B2 => n17380, ZN => n16989);
   U11927 : NOR2_X1 port map( A1 => n16989, A2 => n16597, ZN => DataMem_N1693);
   U11883 : NOR2_X1 port map( A1 => n16989, A2 => n16596, ZN => DataMem_N1757);
   U11848 : NOR2_X1 port map( A1 => n16989, A2 => n16595, ZN => DataMem_N1821);
   U11813 : NOR2_X1 port map( A1 => n16989, A2 => n16594, ZN => DataMem_N1885);
   U11929 : NOR2_X1 port map( A1 => n16990, A2 => n16597, ZN => DataMem_N1691);
   U11779 : NOR2_X1 port map( A1 => n16989, A2 => n16593, ZN => DataMem_N1949);
   U11744 : NOR2_X1 port map( A1 => n16989, A2 => n16592, ZN => DataMem_N2013);
   U11714 : NOR2_X1 port map( A1 => n16994, A2 => n16591, ZN => DataMem_N2067);
   U11709 : NOR2_X1 port map( A1 => n16989, A2 => n16591, ZN => DataMem_N2077);
   U11675 : NOR2_X1 port map( A1 => n16989, A2 => n16590, ZN => DataMem_N2141);
   U11784 : NOR2_X1 port map( A1 => n16994, A2 => n16593, ZN => DataMem_N1939);
   U11539 : AOI22_X1 port map( A1 => n17660, A2 => DataMem_Mem_7_21_port, B1 =>
                           n17530, B2 => DataMem_Mem_6_21_port, ZN => n16871);
   U11538 : AOI22_X1 port map( A1 => n16821, A2 => DataMem_Mem_5_21_port, B1 =>
                           n16822, B2 => DataMem_Mem_4_21_port, ZN => n16872);
   U11537 : AOI22_X1 port map( A1 => n17122, A2 => DataMem_Mem_3_21_port, B1 =>
                           n16820, B2 => DataMem_Mem_2_21_port, ZN => n16873);
   U11536 : AOI22_X1 port map( A1 => n17124, A2 => DataMem_Mem_1_21_port, B1 =>
                           n17125, B2 => DataMem_Mem_0_21_port, ZN => n16874);
   U11534 : NOR2_X1 port map( A1 => n17155, A2 => n16870, ZN => DataMem_N2224);
   U11745 : NOR2_X1 port map( A1 => n16990, A2 => n16592, ZN => DataMem_N2011);
   U11884 : NOR2_X1 port map( A1 => n16990, A2 => n16596, ZN => DataMem_N1755);
   U11749 : NOR2_X1 port map( A1 => n16994, A2 => n16592, ZN => DataMem_N2003);
   U11849 : NOR2_X1 port map( A1 => n16990, A2 => n16595, ZN => DataMem_N1819);
   U11814 : NOR2_X1 port map( A1 => n16990, A2 => n16594, ZN => DataMem_N1883);
   U11780 : NOR2_X1 port map( A1 => n16990, A2 => n16593, ZN => DataMem_N1947);
   U8522 : NAND2_X1 port map( A1 => pipeline_MEM_controls_in_MEM_1_port, A2 => 
                           n14105, ZN => n14104);
   U8510 : OAI22_X1 port map( A1 => n14103, A2 => n14104, B1 => n14092, B2 => 
                           n14105, ZN => n14102);
   U8509 : OAI211_X1 port map( C1 => pipeline_WB_controls_in_MEMWB_1_port, C2 
                           => n14093, A => n14090, B => n14102, ZN => 
                           pipeline_cu_hazard_N39);
   U8457 : NOR2_X1 port map( A1 => pipeline_inst_IFID_DEC_30_port, A2 => n14011
                           , ZN => n14008);
   U8456 : NOR4_X1 port map( A1 => n14007, A2 => n14008, A3 => n14009, A4 => 
                           n14010, ZN => n14003);
   U8454 : NAND2_X1 port map( A1 => n14005, A2 => n13989, ZN => n14004);
   U8453 : NAND4_X1 port map( A1 => n14002, A2 => n14003, A3 => n17704, A4 => 
                           n14004, ZN => pipeline_cu_pipeline_N109);
   U8445 : AOI21_X1 port map( B1 => n13980, B2 => n13984, A => Rst, ZN => 
                           pipeline_cu_pipeline_N113);
   U8443 : NAND2_X1 port map( A1 => n13982, A2 => n13983, ZN => 
                           pipeline_cu_pipeline_N112);
   U10220 : NOR3_X1 port map( A1 => n17347, A2 => n17313, A3 => n14177, ZN => 
                           n14127);
   U10231 : NOR2_X1 port map( A1 => pipeline_stall, A2 => n15648, ZN => n15601)
                           ;
   U11463 : NOR2_X1 port map( A1 => pipeline_RegDst_to_WB_3_port, A2 => 
                           pipeline_RegDst_to_WB_4_port, ZN => n16584);
   U8654 : NOR2_X1 port map( A1 => pipeline_inst_IFID_DEC_29_port, A2 => n14169
                           , ZN => n14007);
   U8633 : NOR4_X1 port map( A1 => n14007, A2 => n14009, A3 => n14183, A4 => 
                           n14184, ZN => n13980);
   U8615 : NOR3_X1 port map( A1 => pipeline_inst_IFID_DEC_27_port, A2 => n14176
                           , A3 => n14177, ZN => pipeline_cu_pipeline_N89);
   U9475 : NAND2_X1 port map( A1 => n17703, A2 => 
                           pipeline_WB_controls_in_MEMWB_1_port, ZN => n14129);
   U11950 : AOI22_X1 port map( A1 => n17744, A2 => 
                           pipeline_data_to_RF_from_WB_11_port, B1 => n13818, 
                           B2 => n17743, ZN => n17000);
   U11952 : AOI22_X1 port map( A1 => pipeline_Forward_sw1_mux, A2 => 
                           pipeline_data_to_RF_from_WB_10_port, B1 => n13816, 
                           B2 => n17743, ZN => n17001);
   U11948 : AOI22_X1 port map( A1 => pipeline_Forward_sw1_mux, A2 => 
                           pipeline_data_to_RF_from_WB_12_port, B1 => n13812, 
                           B2 => n17380, ZN => n16999);
   U11968 : AOI22_X1 port map( A1 => n17744, A2 => 
                           pipeline_data_to_RF_from_WB_2_port, B1 => n13808, B2
                           => n17743, ZN => n17009);
   U11966 : AOI22_X1 port map( A1 => n17744, A2 => 
                           pipeline_data_to_RF_from_WB_3_port, B1 => n13807, B2
                           => n17743, ZN => n17008);
   U11970 : AOI22_X1 port map( A1 => pipeline_Forward_sw1_mux, A2 => 
                           pipeline_data_to_RF_from_WB_1_port, B1 => n13805, B2
                           => n17743, ZN => n17010);
   U11958 : AOI22_X1 port map( A1 => n17744, A2 => 
                           pipeline_data_to_RF_from_WB_7_port, B1 => n13830, B2
                           => n17743, ZN => n17004);
   U11964 : AOI22_X1 port map( A1 => n17744, A2 => 
                           pipeline_data_to_RF_from_WB_4_port, B1 => n13835, B2
                           => n17743, ZN => n17007);
   U11960 : AOI22_X1 port map( A1 => n17744, A2 => 
                           pipeline_data_to_RF_from_WB_6_port, B1 => n13828, B2
                           => n17743, ZN => n17005);
   U11962 : AOI22_X1 port map( A1 => n17744, A2 => 
                           pipeline_data_to_RF_from_WB_5_port, B1 => n13831, B2
                           => n17743, ZN => n17006);
   U11954 : AOI22_X1 port map( A1 => pipeline_Forward_sw1_mux, A2 => 
                           pipeline_data_to_RF_from_WB_9_port, B1 => n13819, B2
                           => n17743, ZN => n17002);
   U11912 : AOI22_X1 port map( A1 => n17744, A2 => 
                           pipeline_data_to_RF_from_WB_30_port, B1 => n13791, 
                           B2 => n17380, ZN => n16981);
   U11956 : AOI22_X1 port map( A1 => n17744, A2 => 
                           pipeline_data_to_RF_from_WB_8_port, B1 => n13785, B2
                           => n17743, ZN => n17003);
   U11914 : AOI22_X1 port map( A1 => pipeline_Forward_sw1_mux, A2 => 
                           pipeline_data_to_RF_from_WB_29_port, B1 => n13792, 
                           B2 => n17743, ZN => n16982);
   U11976 : AOI22_X1 port map( A1 => n17744, A2 => 
                           pipeline_data_to_RF_from_WB_0_port, B1 => n13784, B2
                           => n17743, ZN => n17011);
   U11922 : AOI22_X1 port map( A1 => n17744, A2 => 
                           pipeline_data_to_RF_from_WB_25_port, B1 => n13795, 
                           B2 => n17743, ZN => n16986);
   U11916 : AOI22_X1 port map( A1 => n17744, A2 => 
                           pipeline_data_to_RF_from_WB_28_port, B1 => n13787, 
                           B2 => n17380, ZN => n16983);
   U11924 : AOI22_X1 port map( A1 => n17744, A2 => 
                           pipeline_data_to_RF_from_WB_24_port, B1 => n13786, 
                           B2 => n17743, ZN => n16987);
   U11944 : AOI22_X1 port map( A1 => n17744, A2 => 
                           pipeline_data_to_RF_from_WB_14_port, B1 => n13788, 
                           B2 => n17380, ZN => n16997);
   U11942 : AOI22_X1 port map( A1 => pipeline_Forward_sw1_mux, A2 => 
                           pipeline_data_to_RF_from_WB_15_port, B1 => n13789, 
                           B2 => n17380, ZN => n16996);
   U11930 : AOI22_X1 port map( A1 => n17744, A2 => 
                           pipeline_data_to_RF_from_WB_21_port, B1 => n13798, 
                           B2 => n17380, ZN => n16990);
   U11938 : AOI22_X1 port map( A1 => pipeline_Forward_sw1_mux, A2 => 
                           pipeline_data_to_RF_from_WB_17_port, B1 => n13802, 
                           B2 => n17380, ZN => n16994);
   U11932 : AOI22_X1 port map( A1 => n17744, A2 => 
                           pipeline_data_to_RF_from_WB_20_port, B1 => n13799, 
                           B2 => n17380, ZN => n16991);
   U11926 : AOI22_X1 port map( A1 => n17744, A2 => 
                           pipeline_data_to_RF_from_WB_23_port, B1 => n13796, 
                           B2 => n17743, ZN => n16988);
   U12241 : NAND3_X1 port map( A1 => pipeline_RegDst_to_WB_3_port, A2 => 
                           pipeline_RegDst_to_WB_4_port, A3 => n17643, ZN => 
                           n16589);
   U12234 : NAND3_X1 port map( A1 => pipeline_RegDst_to_WB_4_port, A2 => n17643
                           , A3 => n17385, ZN => n16588);
   U12233 : NAND3_X1 port map( A1 => pipeline_RegDst_to_WB_3_port, A2 => n17643
                           , A3 => n17386, ZN => n16587);
   U10247 : NOR2_X1 port map( A1 => pipeline_inst_IFID_DEC_31_port, A2 => 
                           n17348, ZN => n14049);
   U10244 : NOR2_X1 port map( A1 => n14186, A2 => n14059, ZN => n14126);
   U10240 : NOR2_X1 port map( A1 => pipeline_inst_IFID_DEC_30_port, A2 => 
                           pipeline_inst_IFID_DEC_26_port, ZN => n13993);
   U9893 : NOR2_X1 port map( A1 => Rst, A2 => 
                           pipeline_EXE_controls_in_EXEcute_5_port, ZN => 
                           n14995);
   U9871 : NAND2_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_2_port, A2
                           => n15573, ZN => n14981);
   U9389 : NAND2_X1 port map( A1 => 
                           pipeline_stageD_offset_jump_sign_ext_18_port, A2 => 
                           pipeline_stageD_offset_jump_sign_ext_17_port, ZN => 
                           n14863);
   U9383 : NAND2_X1 port map( A1 => 
                           pipeline_stageD_offset_jump_sign_ext_18_port, A2 => 
                           n17329, ZN => n14865);
   U9371 : NAND2_X1 port map( A1 => 
                           pipeline_stageD_offset_jump_sign_ext_17_port, A2 => 
                           n17408, ZN => n14864);
   U11426 : NOR2_X1 port map( A1 => n16785, A2 => n16786, ZN => n16778);
   U10212 : NOR2_X1 port map( A1 => n15827, A2 => n15828, ZN => n15606);
   U11978 : NAND3_X1 port map( A1 => 
                           pipeline_stageD_offset_to_jump_temp_15_port, A2 => 
                           pipeline_EXE_controls_in_IDEX_8_port, A3 => n13967, 
                           ZN => n13969);
   U8431 : OAI21_X1 port map( B1 => n13967, B2 => n17328, A => n13969, ZN => 
                           pipeline_stageD_offset_to_jump_temp_30_port);
   U10922 : NAND2_X1 port map( A1 => pipeline_WB_controls_in_MEMWB_1_port, A2 
                           => n14103, ZN => n15827);
   U10237 : OAI21_X1 port map( B1 => n15839, B2 => n15840, A => n15841, ZN => 
                           n15838);
   U10213 : NOR2_X1 port map( A1 => n15829, A2 => n15828, ZN => n15605);
   U10902 : NOR2_X1 port map( A1 => n16546, A2 => n16532, ZN => n15930);
   U10901 : NOR2_X1 port map( A1 => n16545, A2 => n16532, ZN => n15931);
   U10899 : NOR2_X1 port map( A1 => n16530, A2 => n16540, ZN => n15928);
   U10898 : NOR2_X1 port map( A1 => n16530, A2 => n16539, ZN => n15929);
   U10896 : NOR2_X1 port map( A1 => n16529, A2 => n16540, ZN => n15926);
   U10895 : NOR2_X1 port map( A1 => n16529, A2 => n16539, ZN => n15927);
   U10893 : NOR2_X1 port map( A1 => n16532, A2 => n16540, ZN => n15924);
   U10892 : NOR2_X1 port map( A1 => n16532, A2 => n16539, ZN => n15925);
   U10929 : NOR4_X1 port map( A1 => n16560, A2 => n16561, A3 => n16562, A4 => 
                           n16563, ZN => n15830);
   U10915 : NOR2_X1 port map( A1 => n16546, A2 => n16530, ZN => n15940);
   U10914 : NOR2_X1 port map( A1 => n16530, A2 => n16545, ZN => n15941);
   U10912 : NAND2_X1 port map( A1 => 
                           pipeline_stageD_offset_jump_sign_ext_23_port, A2 => 
                           n17317, ZN => n16529);
   U10911 : NOR2_X1 port map( A1 => n16546, A2 => n16529, ZN => n15938);
   U10910 : NOR2_X1 port map( A1 => n16545, A2 => n16529, ZN => n15939);
   U10889 : NOR2_X1 port map( A1 => n16527, A2 => n16540, ZN => n15918);
   U10885 : NOR2_X1 port map( A1 => n16532, A2 => n16531, ZN => n15917);
   U10883 : NOR2_X1 port map( A1 => n16533, A2 => n16529, ZN => n15914);
   U10880 : NOR2_X1 port map( A1 => n16533, A2 => n16530, ZN => n15912);
   U10249 : OAI21_X1 port map( B1 => n15830, B2 => n15842, A => n15843, ZN => 
                           n15839);
   U10916 : NAND2_X1 port map( A1 => 
                           pipeline_stageD_offset_jump_sign_ext_22_port, A2 => 
                           pipeline_stageD_offset_jump_sign_ext_23_port, ZN => 
                           n16530);
   U10908 : NAND2_X1 port map( A1 => n17317, A2 => n17383, ZN => n16527);
   U10907 : NOR2_X1 port map( A1 => n16527, A2 => n16533, ZN => n15935);
   U10906 : NOR2_X1 port map( A1 => n16527, A2 => n16546, ZN => n15936);
   U10905 : NOR2_X1 port map( A1 => n16527, A2 => n16545, ZN => n15937);
   U10903 : NAND2_X1 port map( A1 => 
                           pipeline_stageD_offset_jump_sign_ext_22_port, A2 => 
                           n17383, ZN => n16532);
   U10876 : NOR2_X1 port map( A1 => n16529, A2 => n16534, ZN => n15906);
   U10872 : NOR2_X1 port map( A1 => n16532, A2 => n16528, ZN => n15905);
   U10869 : NOR2_X1 port map( A1 => n16530, A2 => n16528, ZN => n15903);
   U10233 : OAI21_X1 port map( B1 => n15834, B2 => n14947, A => n17703, ZN => 
                           n15648);
   U10236 : AOI21_X1 port map( B1 => n13979, B2 => n15646, A => n15838, ZN => 
                           n15834);
   U8441 : INV_X1 port map( A => n13979, ZN => n13967);
   U10936 : INV_X1 port map( A => n16555, ZN => n16560);
   U10766 : INV_X1 port map( A => n15827, ZN => n15832);
   U10746 : INV_X1 port map( A => n14945, ZN => n15772);
   U10726 : INV_X1 port map( A => n14883, ZN => n15688);
   U10260 : INV_X1 port map( A => n15886, ZN => n15842);
   U10239 : INV_X1 port map( A => n13993, ZN => n14176);
   U10224 : INV_X1 port map( A => n15834, ZN => n15833);
   U10218 : NAND2_X1 port map( A1 => n15833, A2 => n14127, ZN => n15828);
   U10214 : INV_X1 port map( A => n15830, ZN => n15829);
   U11317 : INV_X1 port map( A => n15427, ZN => n15426);
   U11313 : OAI21_X1 port map( B1 => n17662, B2 => n17344, A => n16729, ZN => 
                           pipeline_stageE_input1_to_ALU_13_port);
   U11218 : INV_X1 port map( A => pipeline_stageE_input1_to_ALU_4_port, ZN => 
                           n15564);
   U11217 : OR2_X1 port map( A1 => n16683, A2 => n15564, ZN => n15569);
   U11209 : INV_X1 port map( A => n15538, ZN => n15537);
   U11201 : OR2_X1 port map( A1 => pipeline_stageE_input1_to_ALU_6_port, A2 => 
                           n16676, ZN => n15527);
   U11289 : INV_X1 port map( A => n15498, ZN => n15505);
   U11287 : OR2_X1 port map( A1 => pipeline_stageE_input1_to_ALU_8_port, A2 => 
                           n16672, ZN => n15509);
   U11187 : INV_X1 port map( A => n15492, ZN => n15491);
   U11184 : INV_X1 port map( A => n15477, ZN => n15495);
   U11174 : INV_X1 port map( A => n15435, ZN => n15442);
   U11167 : INV_X1 port map( A => n15431, ZN => n15446);
   U11164 : INV_X1 port map( A => n15414, ZN => n15432);
   U11158 : INV_X1 port map( A => n15411, ZN => n15410);
   U11151 : INV_X1 port map( A => n15400, ZN => n15413);
   U11134 : INV_X1 port map( A => n15363, ZN => n15362);
   U11131 : INV_X1 port map( A => n16632, ZN => n15367);
   U11123 : INV_X1 port map( A => n15372, ZN => n15379);
   U11121 : OR2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_A_16_port, A2 
                           => n15369, ZN => n15383);
   U11111 : INV_X1 port map( A => n15331, ZN => n15330);
   U11335 : OAI21_X1 port map( B1 => n17105, B2 => n17322, A => n16738, ZN => 
                           pipeline_stageE_input1_to_ALU_20_port);
   U11353 : INV_X1 port map( A => n15279, ZN => n15278);
   U11089 : OAI21_X1 port map( B1 => n17662, B2 => n17324, A => n16618, ZN => 
                           pipeline_stageE_input1_to_ALU_24_port);
   U11083 : INV_X1 port map( A => n15246, ZN => n15245);
   U11081 : INV_X1 port map( A => n15249, ZN => n16613);
   U11368 : OAI21_X1 port map( B1 => n17662, B2 => n17427, A => n16754, ZN => 
                           pipeline_stageE_input1_to_ALU_25_port);
   U11390 : OR2_X1 port map( A1 => n16611, A2 => 
                           pipeline_stageE_input1_to_ALU_28_port, ZN => n15166)
                           ;
   U9653 : INV_X1 port map( A => n15221, ZN => n15219);
   U9703 : INV_X1 port map( A => n15301, ZN => n15300);
   U9806 : INV_X1 port map( A => n15476, ZN => n15462);
   U9859 : INV_X1 port map( A => n15540, ZN => n15555);
   U9897 : INV_X1 port map( A => n15056, ZN => n15594);
   U9511 : INV_X1 port map( A => n15055, ZN => n15054);
   U9717 : INV_X1 port map( A => n15297, ZN => n15320);
   U11403 : INV_X1 port map( A => n15169, ZN => n15176);
   U9611 : INV_X1 port map( A => n15162, ZN => n15145);
   U11411 : INV_X1 port map( A => n15150, ZN => n15157);
   U11063 : INV_X1 port map( A => n15134, ZN => n15133);
   U10052 : INV_X1 port map( A => n14889, ZN => n15692);
   U10058 : INV_X1 port map( A => n14891, ZN => n15697);
   U9889 : INV_X1 port map( A => n15588, ZN => n15573);
   U9867 : INV_X1 port map( A => n14949, ZN => n14993);
   U10064 : INV_X1 port map( A => n14893, ZN => n15702);
   U9630 : INV_X1 port map( A => n15182, ZN => n15189);
   U10070 : INV_X1 port map( A => n14895, ZN => n15707);
   U9640 : INV_X1 port map( A => n15202, ZN => n15201);
   U9650 : INV_X1 port map( A => n15216, ZN => n15215);
   U10076 : INV_X1 port map( A => n14897, ZN => n15712);
   U9677 : INV_X1 port map( A => n15261, ZN => n15260);
   U9659 : INV_X1 port map( A => n15224, ZN => n15231);
   U10082 : INV_X1 port map( A => n14899, ZN => n15717);
   U9711 : INV_X1 port map( A => n15312, ZN => n15311);
   U9699 : INV_X1 port map( A => n15285, ZN => n15292);
   U9792 : INV_X1 port map( A => n15449, ZN => n15456);
   U9732 : INV_X1 port map( A => n15346, ZN => n15345);
   U9776 : INV_X1 port map( A => pipeline_stageE_input1_to_ALU_13_port, ZN => 
                           n15425);
   U9759 : INV_X1 port map( A => n15386, ZN => n15393);
   U10088 : INV_X1 port map( A => n14901, ZN => n15722);
   U9856 : INV_X1 port map( A => n15553, ZN => n15552);
   U9805 : INV_X1 port map( A => n15474, ZN => n15473);
   U9832 : INV_X1 port map( A => n15512, ZN => n15519);
   U10094 : INV_X1 port map( A => n14903, ZN => n15727);
   U9980 : INV_X1 port map( A => n15653, ZN => n3957);
   U9972 : INV_X1 port map( A => n15649, ZN => n3961);
   U9968 : INV_X1 port map( A => n15645, ZN => n3963);
   U9960 : INV_X1 port map( A => n15641, ZN => n3967);
   U9976 : INV_X1 port map( A => n15651, ZN => n3959);
   U9962 : INV_X1 port map( A => n15642, ZN => n3966);
   U10144 : INV_X1 port map( A => n15768, ZN => n3881);
   U10155 : INV_X1 port map( A => n15778, ZN => n3877);
   U10066 : INV_X1 port map( A => n15703, ZN => n3907);
   U9940 : INV_X1 port map( A => n15631, ZN => n3977);
   U9964 : INV_X1 port map( A => n15643, ZN => n3965);
   U10054 : INV_X1 port map( A => n15693, ZN => n3911);
   U10197 : INV_X1 port map( A => n15813, ZN => n3863);
   U10173 : INV_X1 port map( A => n15793, ZN => n3871);
   U9930 : INV_X1 port map( A => n15626, ZN => n3982);
   U10090 : INV_X1 port map( A => n15723, ZN => n3899);
   U10108 : INV_X1 port map( A => n15738, ZN => n3893);
   U9952 : INV_X1 port map( A => n15637, ZN => n3971);
   U10167 : INV_X1 port map( A => n15788, ZN => n3873);
   U9928 : INV_X1 port map( A => n15625, ZN => n3983);
   U10078 : INV_X1 port map( A => n15713, ZN => n3903);
   U10138 : INV_X1 port map( A => n15763, ZN => n3883);
   U9904 : INV_X1 port map( A => n15599, ZN => n3992);
   U9950 : INV_X1 port map( A => n15636, ZN => n3972);
   U10161 : INV_X1 port map( A => n15783, ZN => n3875);
   U10229 : INV_X1 port map( A => n15837, ZN => n3855);
   U9956 : INV_X1 port map( A => n15639, ZN => n3969);
   U10209 : INV_X1 port map( A => n15823, ZN => n3859);
   U9958 : INV_X1 port map( A => n15640, ZN => n3968);
   U10126 : INV_X1 port map( A => n15753, ZN => n3887);
   U10120 : INV_X1 port map( A => n15748, ZN => n3889);
   U10102 : INV_X1 port map( A => n15733, ZN => n3895);
   U9938 : INV_X1 port map( A => n15630, ZN => n3978);
   U9946 : INV_X1 port map( A => n15634, ZN => n3974);
   U9942 : INV_X1 port map( A => n15632, ZN => n3976);
   U10072 : INV_X1 port map( A => n15708, ZN => n3905);
   U10096 : INV_X1 port map( A => n15728, ZN => n3897);
   U9922 : INV_X1 port map( A => n15622, ZN => n3986);
   U9932 : INV_X1 port map( A => n15627, ZN => n3981);
   U9944 : INV_X1 port map( A => n15633, ZN => n3975);
   U10060 : INV_X1 port map( A => n15698, ZN => n3909);
   U10203 : INV_X1 port map( A => n15818, ZN => n3861);
   U10191 : INV_X1 port map( A => n15808, ZN => n3865);
   U10185 : INV_X1 port map( A => n15803, ZN => n3867);
   U10225 : INV_X1 port map( A => n15835, ZN => n3857);
   U10149 : INV_X1 port map( A => n15773, ZN => n3879);
   U9924 : INV_X1 port map( A => n15623, ZN => n3985);
   U9954 : INV_X1 port map( A => n15638, ZN => n3970);
   U9948 : INV_X1 port map( A => n15635, ZN => n3973);
   U10100 : INV_X1 port map( A => n14905, ZN => n15732);
   U10049 : AND2_X1 port map( A1 => n15600, A2 => n13937, ZN => n3923);
   U10201 : INV_X1 port map( A => n14921, ZN => n15817);
   U10142 : INV_X1 port map( A => n14929, ZN => n15767);
   U10112 : INV_X1 port map( A => n14909, ZN => n15742);
   U10124 : INV_X1 port map( A => n14915, ZN => n15752);
   U10153 : INV_X1 port map( A => n14939, ZN => n15777);
   U9908 : INV_X1 port map( A => n14913, ZN => n15609);
   U10195 : INV_X1 port map( A => n14925, ZN => n15812);
   U10165 : INV_X1 port map( A => n14937, ZN => n15787);
   U10207 : INV_X1 port map( A => n14941, ZN => n15822);
   U10132 : INV_X1 port map( A => n15758, ZN => n3885);
   U10114 : INV_X1 port map( A => n15743, ZN => n3891);
   U9936 : INV_X1 port map( A => n15629, ZN => n3979);
   U10227 : INV_X1 port map( A => n15836, ZN => n3856);
   U10177 : INV_X1 port map( A => n14933, ZN => n15797);
   U10136 : INV_X1 port map( A => n14919, ZN => n15762);
   U10106 : INV_X1 port map( A => n14907, ZN => n15737);
   U10171 : INV_X1 port map( A => n14935, ZN => n15792);
   U10159 : INV_X1 port map( A => n14931, ZN => n15782);
   U10118 : INV_X1 port map( A => n14911, ZN => n15747);
   U10216 : INV_X1 port map( A => n14943, ZN => n15831);
   U10183 : INV_X1 port map( A => n14923, ZN => n15802);
   U10130 : INV_X1 port map( A => n14917, ZN => n15757);
   U10189 : INV_X1 port map( A => n14927, ZN => n15807);
   U9966 : INV_X1 port map( A => n15644, ZN => n3964);
   U9934 : INV_X1 port map( A => n15628, ZN => n3980);
   U9926 : INV_X1 port map( A => n15624, ZN => n3984);
   U9910 : INV_X1 port map( A => n15612, ZN => n3990);
   U10179 : INV_X1 port map( A => n15798, ZN => n3869);
   U10084 : INV_X1 port map( A => n15718, ZN => n3901);
   U9456 : INV_X1 port map( A => n14947, ZN => n14025);
   U8652 : INV_X1 port map( A => n13998, ZN => n14001);
   U8646 : INV_X1 port map( A => n14011, ZN => n14185);
   U8623 : AND2_X1 port map( A1 => n17412, A2 => n14179, ZN => n14044);
   U8593 : INV_X1 port map( A => n14165, ZN => pipeline_MEMWB_Stage_N12);
   U8595 : INV_X1 port map( A => n14166, ZN => pipeline_MEMWB_Stage_N11);
   U8565 : INV_X1 port map( A => n14151, ZN => pipeline_MEMWB_Stage_N26);
   U8569 : INV_X1 port map( A => n14153, ZN => pipeline_MEMWB_Stage_N24);
   U8547 : INV_X1 port map( A => n14142, ZN => pipeline_MEMWB_Stage_N35);
   U8583 : INV_X1 port map( A => n14160, ZN => pipeline_MEMWB_Stage_N17);
   U8539 : INV_X1 port map( A => n14138, ZN => pipeline_MEMWB_Stage_N39);
   U8571 : INV_X1 port map( A => n14154, ZN => pipeline_MEMWB_Stage_N23);
   U8533 : INV_X1 port map( A => n14133, ZN => pipeline_MEMWB_Stage_N42);
   U8545 : INV_X1 port map( A => n14141, ZN => pipeline_MEMWB_Stage_N36);
   U8549 : INV_X1 port map( A => n14143, ZN => pipeline_MEMWB_Stage_N34);
   U8587 : INV_X1 port map( A => n14162, ZN => pipeline_MEMWB_Stage_N15);
   U8589 : INV_X1 port map( A => n14163, ZN => pipeline_MEMWB_Stage_N14);
   U8579 : INV_X1 port map( A => n14158, ZN => pipeline_MEMWB_Stage_N19);
   U8581 : INV_X1 port map( A => n14159, ZN => pipeline_MEMWB_Stage_N18);
   U8551 : INV_X1 port map( A => n14144, ZN => pipeline_MEMWB_Stage_N33);
   U8591 : INV_X1 port map( A => n14164, ZN => pipeline_MEMWB_Stage_N13);
   U8577 : INV_X1 port map( A => n14157, ZN => pipeline_MEMWB_Stage_N20);
   U8553 : INV_X1 port map( A => n14145, ZN => pipeline_MEMWB_Stage_N32);
   U8573 : INV_X1 port map( A => n14155, ZN => pipeline_MEMWB_Stage_N22);
   U8559 : INV_X1 port map( A => n14148, ZN => pipeline_MEMWB_Stage_N29);
   U8555 : INV_X1 port map( A => n14146, ZN => pipeline_MEMWB_Stage_N31);
   U8535 : INV_X1 port map( A => n14136, ZN => pipeline_MEMWB_Stage_N41);
   U8537 : INV_X1 port map( A => n14137, ZN => pipeline_MEMWB_Stage_N40);
   U8541 : INV_X1 port map( A => n14139, ZN => pipeline_MEMWB_Stage_N38);
   U8557 : INV_X1 port map( A => n14147, ZN => pipeline_MEMWB_Stage_N30);
   U8543 : INV_X1 port map( A => n14140, ZN => pipeline_MEMWB_Stage_N37);
   U8567 : INV_X1 port map( A => n14152, ZN => pipeline_MEMWB_Stage_N25);
   U8585 : INV_X1 port map( A => n14161, ZN => pipeline_MEMWB_Stage_N16);
   U8561 : INV_X1 port map( A => n14149, ZN => pipeline_MEMWB_Stage_N28);
   U8563 : INV_X1 port map( A => n14150, ZN => pipeline_MEMWB_Stage_N27);
   U8575 : INV_X1 port map( A => n14156, ZN => pipeline_MEMWB_Stage_N21);
   U8604 : AND2_X1 port map( A1 => n14167, A2 => 
                           pipeline_EXE_controls_in_IDEX_2_port, ZN => 
                           pipeline_IDEX_Stage_N95);
   U8601 : AND2_X1 port map( A1 => n14167, A2 => 
                           pipeline_EXE_controls_in_IDEX_5_port, ZN => 
                           pipeline_IDEX_Stage_N98);
   U8602 : AND2_X1 port map( A1 => n14167, A2 => 
                           pipeline_EXE_controls_in_IDEX_4_port, ZN => 
                           pipeline_IDEX_Stage_N97);
   U9458 : AND2_X1 port map( A1 => n14167, A2 => 
                           pipeline_EXE_controls_in_IDEX_7_port, ZN => 
                           pipeline_IDEX_Stage_N100);
   U9457 : AND2_X1 port map( A1 => n14167, A2 => 
                           pipeline_EXE_controls_in_IDEX_8_port, ZN => 
                           pipeline_IDEX_Stage_N101);
   U8600 : AND2_X1 port map( A1 => n14167, A2 => 
                           pipeline_EXE_controls_in_IDEX_6_port, ZN => 
                           pipeline_IDEX_Stage_N99);
   U8603 : AND2_X1 port map( A1 => n14167, A2 => 
                           pipeline_EXE_controls_in_IDEX_3_port, ZN => 
                           pipeline_IDEX_Stage_N96);
   U8656 : AND2_X1 port map( A1 => n14167, A2 => 
                           pipeline_WB_controls_in_IDEX_0_port, ZN => 
                           pipeline_IDEX_Stage_N89);
   U8605 : AND2_X1 port map( A1 => n14167, A2 => 
                           pipeline_EXE_controls_in_IDEX_1_port, ZN => 
                           pipeline_IDEX_Stage_N94);
   U8606 : AND2_X1 port map( A1 => n14167, A2 => 
                           pipeline_EXE_controls_in_IDEX_0_port, ZN => 
                           pipeline_IDEX_Stage_N93);
   U8610 : INV_X1 port map( A => n14123, ZN => n13981);
   U8599 : INV_X1 port map( A => n14129, ZN => pipeline_MEMWB_Stage_N10);
   U8532 : AND2_X1 port map( A1 => pipeline_regDst_to_mem_0_port, A2 => 
                           pipeline_MEMWB_Stage_N10, ZN => 
                           pipeline_MEMWB_Stage_N43);
   U9477 : INV_X1 port map( A => n14120, ZN => n14101);
   U9682 : AND2_X1 port map( A1 => n13936, A2 => n17705, ZN => 
                           pipeline_EXMEM_stage_N3);
   U9542 : AND2_X1 port map( A1 => pipeline_MEM_controls_in_EXMEM_1_port, A2 =>
                           n17705, ZN => pipeline_EXMEM_stage_N6);
   U11975 : NOR3_X2 port map( A1 => addr_to_dataRam_4_port, A2 => 
                           addr_to_dataRam_2_port, A3 => addr_to_dataRam_3_port
                           , ZN => n16818);
   U11907 : NOR3_X2 port map( A1 => addr_to_dataRam_4_port, A2 => 
                           addr_to_dataRam_3_port, A3 => n17012, ZN => n16817);
   U11595 : AND4_X1 port map( A1 => n16921, A2 => n16922, A3 => n16923, A4 => 
                           n16924, ZN => n16920);
   U11589 : AND4_X1 port map( A1 => n16916, A2 => n16917, A3 => n16918, A4 => 
                           n16919, ZN => n16915);
   U11649 : AND4_X1 port map( A1 => n16966, A2 => n16967, A3 => n16968, A4 => 
                           n16969, ZN => n16965);
   U11643 : AND4_X1 port map( A1 => n16961, A2 => n16962, A3 => n16963, A4 => 
                           n16964, ZN => n16960);
   U11637 : AND4_X1 port map( A1 => n16956, A2 => n16957, A3 => n16958, A4 => 
                           n16959, ZN => n16955);
   U11601 : AND4_X1 port map( A1 => n16926, A2 => n16927, A3 => n16928, A4 => 
                           n16929, ZN => n16925);
   U11619 : AND4_X1 port map( A1 => n16941, A2 => n16942, A3 => n16943, A4 => 
                           n16944, ZN => n16940);
   U11631 : AND4_X1 port map( A1 => n16951, A2 => n16952, A3 => n16953, A4 => 
                           n16954, ZN => n16950);
   U11607 : AND4_X1 port map( A1 => n16931, A2 => n16932, A3 => n16933, A4 => 
                           n16934, ZN => n16930);
   U11655 : AND4_X1 port map( A1 => n16971, A2 => n16972, A3 => n16973, A4 => 
                           n16974, ZN => n16970);
   U11625 : AND4_X1 port map( A1 => n16946, A2 => n16947, A3 => n16948, A4 => 
                           n16949, ZN => n16945);
   U11487 : AND4_X1 port map( A1 => n16831, A2 => n16832, A3 => n16833, A4 => 
                           n16834, ZN => n16830);
   U11613 : AND4_X1 port map( A1 => n16936, A2 => n16937, A3 => n16938, A4 => 
                           n16939, ZN => n16935);
   U11499 : AND4_X1 port map( A1 => n16841, A2 => n16842, A3 => n16843, A4 => 
                           n16844, ZN => n16840);
   U11505 : AND4_X1 port map( A1 => n16846, A2 => n16847, A3 => n16848, A4 => 
                           n16849, ZN => n16845);
   U11661 : AND4_X1 port map( A1 => n16976, A2 => n16977, A3 => n16978, A4 => 
                           n16979, ZN => n16975);
   U11511 : AND4_X1 port map( A1 => n16851, A2 => n16852, A3 => n16853, A4 => 
                           n16854, ZN => n16850);
   U11577 : AND4_X1 port map( A1 => n16906, A2 => n16907, A3 => n16908, A4 => 
                           n16909, ZN => n16905);
   U11571 : AND4_X1 port map( A1 => n16901, A2 => n16902, A3 => n16903, A4 => 
                           n16904, ZN => n16900);
   U11517 : AND4_X1 port map( A1 => n16856, A2 => n16857, A3 => n16858, A4 => 
                           n16859, ZN => n16855);
   U11583 : AND4_X1 port map( A1 => n16911, A2 => n16912, A3 => n16913, A4 => 
                           n16914, ZN => n16910);
   U11481 : AND4_X1 port map( A1 => n16826, A2 => n16827, A3 => n16828, A4 => 
                           n16829, ZN => n16825);
   U11493 : AND4_X1 port map( A1 => n16836, A2 => n16837, A3 => n16838, A4 => 
                           n16839, ZN => n16835);
   U11541 : AND4_X1 port map( A1 => n16876, A2 => n16877, A3 => n16878, A4 => 
                           n16879, ZN => n16875);
   U11547 : AND4_X1 port map( A1 => n16881, A2 => n16882, A3 => n16883, A4 => 
                           n16884, ZN => n16880);
   U11559 : AND4_X1 port map( A1 => n16891, A2 => n16892, A3 => n16893, A4 => 
                           n16894, ZN => n16890);
   U8525 : INV_X1 port map( A => n14094, ZN => n14091);
   U8485 : AND3_X1 port map( A1 => n14005, A2 => n14067, A3 => n17350, ZN => 
                           n14033);
   U8466 : AND2_X1 port map( A1 => n13981, A2 => n14030, ZN => n14002);
   U8474 : AND2_X1 port map( A1 => n14051, A2 => n14033, ZN => n14015);
   U8455 : INV_X1 port map( A => n14006, ZN => n13989);
   U8496 : INV_X1 port map( A => pipeline_cu_pipeline_N89, ZN => n13984);
   U11553 : AND4_X1 port map( A1 => n16886, A2 => n16887, A3 => n16888, A4 => 
                           n16889, ZN => n16885);
   U8489 : INV_X1 port map( A => n14005, ZN => n14012);
   U8480 : INV_X1 port map( A => n14061, ZN => n14020);
   U8458 : INV_X1 port map( A => n13988, ZN => pipeline_cu_pipeline_N108);
   U8462 : INV_X1 port map( A => n14022, ZN => n14018);
   U8470 : INV_X1 port map( A => n14040, ZN => n14034);
   U11523 : AND4_X1 port map( A1 => n16861, A2 => n16862, A3 => n16863, A4 => 
                           n16864, ZN => n16860);
   U11475 : AND4_X1 port map( A1 => n16813, A2 => n16814, A3 => n16815, A4 => 
                           n16816, ZN => n16812);
   U11565 : AND4_X1 port map( A1 => n16896, A2 => n16897, A3 => n16898, A4 => 
                           n16899, ZN => n16895);
   U11529 : AND4_X1 port map( A1 => n16866, A2 => n16867, A3 => n16868, A4 => 
                           n16869, ZN => n16865);
   U11535 : AND4_X1 port map( A1 => n16871, A2 => n16872, A3 => n16873, A4 => 
                           n16874, ZN => n16870);
   U8523 : INV_X1 port map( A => n14093, ZN => n14105);
   U8444 : INV_X1 port map( A => pipeline_cu_pipeline_N113, ZN => n13982);
   pipeline_IFID_stage_Instr_out_IFID_reg_0_inst : DFF_X2 port map( D => n3987,
                           CK => Clk, Q => net175543, QN => n17076);
   pipeline_stageF_PC_plus4_add_26_U56 : INV_X1 port map( A => 
                           addr_to_iram_2_port, ZN => 
                           pipeline_stageF_PC_plus4_N9);
   pipeline_stageF_PC_plus4_add_26_U54 : AND2_X1 port map( A1 => 
                           pipeline_stageF_PC_plus4_add_26_carry_28_port, A2 =>
                           addr_to_iram_28_port, ZN => 
                           pipeline_stageF_PC_plus4_add_26_carry_29_port);
   pipeline_stageF_PC_plus4_add_26_U52 : AND2_X1 port map( A1 => 
                           pipeline_stageF_PC_plus4_add_26_carry_27_port, A2 =>
                           addr_to_iram_27_port, ZN => 
                           pipeline_stageF_PC_plus4_add_26_carry_28_port);
   pipeline_stageF_PC_plus4_add_26_U50 : AND2_X1 port map( A1 => 
                           pipeline_stageF_PC_plus4_add_26_carry_26_port, A2 =>
                           addr_to_iram_26_port, ZN => 
                           pipeline_stageF_PC_plus4_add_26_carry_27_port);
   pipeline_stageF_PC_plus4_add_26_U48 : AND2_X1 port map( A1 => 
                           pipeline_stageF_PC_plus4_add_26_carry_25_port, A2 =>
                           addr_to_iram_25_port, ZN => 
                           pipeline_stageF_PC_plus4_add_26_carry_26_port);
   pipeline_stageF_PC_plus4_add_26_U46 : AND2_X1 port map( A1 => 
                           pipeline_stageF_PC_plus4_add_26_carry_24_port, A2 =>
                           addr_to_iram_24_port, ZN => 
                           pipeline_stageF_PC_plus4_add_26_carry_25_port);
   pipeline_stageF_PC_plus4_add_26_U44 : AND2_X1 port map( A1 => 
                           pipeline_stageF_PC_plus4_add_26_carry_23_port, A2 =>
                           addr_to_iram_23_port, ZN => 
                           pipeline_stageF_PC_plus4_add_26_carry_24_port);
   pipeline_stageF_PC_plus4_add_26_U42 : AND2_X1 port map( A1 => 
                           pipeline_stageF_PC_plus4_add_26_carry_22_port, A2 =>
                           addr_to_iram_22_port, ZN => 
                           pipeline_stageF_PC_plus4_add_26_carry_23_port);
   pipeline_stageF_PC_plus4_add_26_U40 : AND2_X1 port map( A1 => 
                           pipeline_stageF_PC_plus4_add_26_carry_21_port, A2 =>
                           addr_to_iram_21_port, ZN => 
                           pipeline_stageF_PC_plus4_add_26_carry_22_port);
   pipeline_stageF_PC_plus4_add_26_U38 : AND2_X1 port map( A1 => 
                           pipeline_stageF_PC_plus4_add_26_carry_20_port, A2 =>
                           addr_to_iram_20_port, ZN => 
                           pipeline_stageF_PC_plus4_add_26_carry_21_port);
   pipeline_stageF_PC_plus4_add_26_U36 : AND2_X1 port map( A1 => 
                           pipeline_stageF_PC_plus4_add_26_carry_19_port, A2 =>
                           addr_to_iram_19_port, ZN => 
                           pipeline_stageF_PC_plus4_add_26_carry_20_port);
   pipeline_stageF_PC_plus4_add_26_U34 : AND2_X1 port map( A1 => 
                           pipeline_stageF_PC_plus4_add_26_carry_18_port, A2 =>
                           addr_to_iram_18_port, ZN => 
                           pipeline_stageF_PC_plus4_add_26_carry_19_port);
   pipeline_stageF_PC_plus4_add_26_U32 : AND2_X1 port map( A1 => 
                           pipeline_stageF_PC_plus4_add_26_carry_17_port, A2 =>
                           addr_to_iram_17_port, ZN => 
                           pipeline_stageF_PC_plus4_add_26_carry_18_port);
   pipeline_stageF_PC_plus4_add_26_U30 : AND2_X1 port map( A1 => 
                           pipeline_stageF_PC_plus4_add_26_carry_16_port, A2 =>
                           addr_to_iram_16_port, ZN => 
                           pipeline_stageF_PC_plus4_add_26_carry_17_port);
   pipeline_stageF_PC_plus4_add_26_U28 : AND2_X1 port map( A1 => 
                           pipeline_stageF_PC_plus4_add_26_carry_15_port, A2 =>
                           addr_to_iram_15_port, ZN => 
                           pipeline_stageF_PC_plus4_add_26_carry_16_port);
   pipeline_stageF_PC_plus4_add_26_U26 : AND2_X1 port map( A1 => 
                           pipeline_stageF_PC_plus4_add_26_carry_14_port, A2 =>
                           addr_to_iram_14_port, ZN => 
                           pipeline_stageF_PC_plus4_add_26_carry_15_port);
   pipeline_stageF_PC_plus4_add_26_U24 : AND2_X1 port map( A1 => 
                           pipeline_stageF_PC_plus4_add_26_carry_13_port, A2 =>
                           addr_to_iram_13_port, ZN => 
                           pipeline_stageF_PC_plus4_add_26_carry_14_port);
   pipeline_stageF_PC_plus4_add_26_U22 : AND2_X1 port map( A1 => 
                           pipeline_stageF_PC_plus4_add_26_carry_12_port, A2 =>
                           addr_to_iram_12_port, ZN => 
                           pipeline_stageF_PC_plus4_add_26_carry_13_port);
   pipeline_stageF_PC_plus4_add_26_U20 : AND2_X1 port map( A1 => 
                           pipeline_stageF_PC_plus4_add_26_carry_11_port, A2 =>
                           addr_to_iram_11_port, ZN => 
                           pipeline_stageF_PC_plus4_add_26_carry_12_port);
   pipeline_stageF_PC_plus4_add_26_U18 : AND2_X1 port map( A1 => 
                           pipeline_stageF_PC_plus4_add_26_carry_10_port, A2 =>
                           addr_to_iram_10_port, ZN => 
                           pipeline_stageF_PC_plus4_add_26_carry_11_port);
   pipeline_stageF_PC_plus4_add_26_U16 : AND2_X1 port map( A1 => 
                           pipeline_stageF_PC_plus4_add_26_carry_9_port, A2 => 
                           addr_to_iram_9_port, ZN => 
                           pipeline_stageF_PC_plus4_add_26_carry_10_port);
   pipeline_stageF_PC_plus4_add_26_U14 : AND2_X1 port map( A1 => 
                           pipeline_stageF_PC_plus4_add_26_carry_8_port, A2 => 
                           addr_to_iram_8_port, ZN => 
                           pipeline_stageF_PC_plus4_add_26_carry_9_port);
   pipeline_stageF_PC_plus4_add_26_U12 : AND2_X1 port map( A1 => 
                           pipeline_stageF_PC_plus4_add_26_carry_7_port, A2 => 
                           addr_to_iram_7_port, ZN => 
                           pipeline_stageF_PC_plus4_add_26_carry_8_port);
   pipeline_stageF_PC_plus4_add_26_U10 : AND2_X1 port map( A1 => 
                           pipeline_stageF_PC_plus4_add_26_carry_6_port, A2 => 
                           addr_to_iram_6_port, ZN => 
                           pipeline_stageF_PC_plus4_add_26_carry_7_port);
   pipeline_stageF_PC_plus4_add_26_U8 : AND2_X1 port map( A1 => 
                           pipeline_stageF_PC_plus4_add_26_carry_5_port, A2 => 
                           addr_to_iram_5_port, ZN => 
                           pipeline_stageF_PC_plus4_add_26_carry_6_port);
   pipeline_stageF_PC_plus4_add_26_U6 : AND2_X1 port map( A1 => 
                           pipeline_stageF_PC_plus4_add_26_carry_4_port, A2 => 
                           addr_to_iram_4_port, ZN => 
                           pipeline_stageF_PC_plus4_add_26_carry_5_port);
   pipeline_stageF_PC_plus4_add_26_U4 : AND2_X1 port map( A1 => 
                           addr_to_iram_2_port, A2 => addr_to_iram_3_port, ZN 
                           => pipeline_stageF_PC_plus4_add_26_carry_4_port);
   pipeline_stageF_PC_plus4_add_26_U1 : XNOR2_X1 port map( A => 
                           addr_to_iram_30_port, B => 
                           pipeline_stageF_PC_plus4_add_26_n1, ZN => 
                           pipeline_stageF_PC_plus4_N37);
   pipeline_stageF_PC_plus4_add_26_U2 : NAND2_X1 port map( A1 => 
                           pipeline_stageF_PC_plus4_add_26_carry_29_port, A2 =>
                           addr_to_iram_29_port, ZN => 
                           pipeline_stageF_PC_plus4_add_26_n1);
   pipeline_stageF_PC_plus4_add_26_U55 : XOR2_X1 port map( A => 
                           addr_to_iram_3_port, B => addr_to_iram_2_port, Z => 
                           pipeline_stageF_PC_plus4_N10);
   pipeline_stageF_PC_plus4_add_26_U53 : XOR2_X1 port map( A => 
                           addr_to_iram_4_port, B => 
                           pipeline_stageF_PC_plus4_add_26_carry_4_port, Z => 
                           pipeline_stageF_PC_plus4_N11);
   pipeline_stageF_PC_plus4_add_26_U51 : XOR2_X1 port map( A => 
                           addr_to_iram_5_port, B => 
                           pipeline_stageF_PC_plus4_add_26_carry_5_port, Z => 
                           pipeline_stageF_PC_plus4_N12);
   pipeline_stageF_PC_plus4_add_26_U49 : XOR2_X1 port map( A => 
                           addr_to_iram_6_port, B => 
                           pipeline_stageF_PC_plus4_add_26_carry_6_port, Z => 
                           pipeline_stageF_PC_plus4_N13);
   pipeline_stageF_PC_plus4_add_26_U47 : XOR2_X1 port map( A => 
                           addr_to_iram_7_port, B => 
                           pipeline_stageF_PC_plus4_add_26_carry_7_port, Z => 
                           pipeline_stageF_PC_plus4_N14);
   pipeline_stageF_PC_plus4_add_26_U45 : XOR2_X1 port map( A => 
                           addr_to_iram_8_port, B => 
                           pipeline_stageF_PC_plus4_add_26_carry_8_port, Z => 
                           pipeline_stageF_PC_plus4_N15);
   pipeline_stageF_PC_plus4_add_26_U43 : XOR2_X1 port map( A => 
                           addr_to_iram_9_port, B => 
                           pipeline_stageF_PC_plus4_add_26_carry_9_port, Z => 
                           pipeline_stageF_PC_plus4_N16);
   pipeline_stageF_PC_plus4_add_26_U41 : XOR2_X1 port map( A => 
                           addr_to_iram_10_port, B => 
                           pipeline_stageF_PC_plus4_add_26_carry_10_port, Z => 
                           pipeline_stageF_PC_plus4_N17);
   pipeline_stageF_PC_plus4_add_26_U39 : XOR2_X1 port map( A => 
                           addr_to_iram_11_port, B => 
                           pipeline_stageF_PC_plus4_add_26_carry_11_port, Z => 
                           pipeline_stageF_PC_plus4_N18);
   pipeline_stageF_PC_plus4_add_26_U37 : XOR2_X1 port map( A => 
                           addr_to_iram_12_port, B => 
                           pipeline_stageF_PC_plus4_add_26_carry_12_port, Z => 
                           pipeline_stageF_PC_plus4_N19);
   pipeline_stageF_PC_plus4_add_26_U35 : XOR2_X1 port map( A => 
                           addr_to_iram_13_port, B => 
                           pipeline_stageF_PC_plus4_add_26_carry_13_port, Z => 
                           pipeline_stageF_PC_plus4_N20);
   pipeline_stageF_PC_plus4_add_26_U33 : XOR2_X1 port map( A => 
                           addr_to_iram_14_port, B => 
                           pipeline_stageF_PC_plus4_add_26_carry_14_port, Z => 
                           pipeline_stageF_PC_plus4_N21);
   pipeline_stageF_PC_plus4_add_26_U31 : XOR2_X1 port map( A => 
                           addr_to_iram_15_port, B => 
                           pipeline_stageF_PC_plus4_add_26_carry_15_port, Z => 
                           pipeline_stageF_PC_plus4_N22);
   pipeline_stageF_PC_plus4_add_26_U29 : XOR2_X1 port map( A => 
                           addr_to_iram_16_port, B => 
                           pipeline_stageF_PC_plus4_add_26_carry_16_port, Z => 
                           pipeline_stageF_PC_plus4_N23);
   pipeline_stageF_PC_plus4_add_26_U27 : XOR2_X1 port map( A => 
                           addr_to_iram_17_port, B => 
                           pipeline_stageF_PC_plus4_add_26_carry_17_port, Z => 
                           pipeline_stageF_PC_plus4_N24);
   pipeline_stageF_PC_plus4_add_26_U25 : XOR2_X1 port map( A => 
                           addr_to_iram_18_port, B => 
                           pipeline_stageF_PC_plus4_add_26_carry_18_port, Z => 
                           pipeline_stageF_PC_plus4_N25);
   pipeline_stageF_PC_plus4_add_26_U23 : XOR2_X1 port map( A => 
                           addr_to_iram_19_port, B => 
                           pipeline_stageF_PC_plus4_add_26_carry_19_port, Z => 
                           pipeline_stageF_PC_plus4_N26);
   pipeline_stageF_PC_plus4_add_26_U21 : XOR2_X1 port map( A => 
                           addr_to_iram_20_port, B => 
                           pipeline_stageF_PC_plus4_add_26_carry_20_port, Z => 
                           pipeline_stageF_PC_plus4_N27);
   pipeline_stageF_PC_plus4_add_26_U19 : XOR2_X1 port map( A => 
                           addr_to_iram_21_port, B => 
                           pipeline_stageF_PC_plus4_add_26_carry_21_port, Z => 
                           pipeline_stageF_PC_plus4_N28);
   pipeline_stageF_PC_plus4_add_26_U17 : XOR2_X1 port map( A => 
                           addr_to_iram_22_port, B => 
                           pipeline_stageF_PC_plus4_add_26_carry_22_port, Z => 
                           pipeline_stageF_PC_plus4_N29);
   pipeline_stageF_PC_plus4_add_26_U15 : XOR2_X1 port map( A => 
                           addr_to_iram_23_port, B => 
                           pipeline_stageF_PC_plus4_add_26_carry_23_port, Z => 
                           pipeline_stageF_PC_plus4_N30);
   pipeline_stageF_PC_plus4_add_26_U13 : XOR2_X1 port map( A => 
                           addr_to_iram_24_port, B => 
                           pipeline_stageF_PC_plus4_add_26_carry_24_port, Z => 
                           pipeline_stageF_PC_plus4_N31);
   pipeline_stageF_PC_plus4_add_26_U11 : XOR2_X1 port map( A => 
                           addr_to_iram_25_port, B => 
                           pipeline_stageF_PC_plus4_add_26_carry_25_port, Z => 
                           pipeline_stageF_PC_plus4_N32);
   pipeline_stageF_PC_plus4_add_26_U9 : XOR2_X1 port map( A => 
                           addr_to_iram_26_port, B => 
                           pipeline_stageF_PC_plus4_add_26_carry_26_port, Z => 
                           pipeline_stageF_PC_plus4_N33);
   pipeline_stageF_PC_plus4_add_26_U7 : XOR2_X1 port map( A => 
                           addr_to_iram_27_port, B => 
                           pipeline_stageF_PC_plus4_add_26_carry_27_port, Z => 
                           pipeline_stageF_PC_plus4_N34);
   pipeline_stageF_PC_plus4_add_26_U5 : XOR2_X1 port map( A => 
                           addr_to_iram_28_port, B => 
                           pipeline_stageF_PC_plus4_add_26_carry_28_port, Z => 
                           pipeline_stageF_PC_plus4_N35);
   pipeline_stageF_PC_plus4_add_26_U3 : XOR2_X1 port map( A => 
                           addr_to_iram_29_port, B => 
                           pipeline_stageF_PC_plus4_add_26_carry_29_port, Z => 
                           pipeline_stageF_PC_plus4_N36);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U97 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n109, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n108);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U92 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n45, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n23);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U85 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n115, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n30);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U162 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n152, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n151);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U91 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n64, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n29);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U29 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n83, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n82);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U86 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n99, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n9);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U93 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n4, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n35);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U112 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n60, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n114);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U45 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n24, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n112);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U44 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n25, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n111);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U165 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n133, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n132);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U89 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n107, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n106);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U11 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n40, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n8);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U26 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n88, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n87);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U107 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n90, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n89);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U104 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n102, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n101);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U111 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n103, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n75);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U94 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n14, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n39);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U12 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n5, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n43);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U87 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n134, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n17);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U168 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n162, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n161);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U95 : AND2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_3_port, A2 
                           => n17302, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n158);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U100 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n164, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n163);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U110 : AND2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_3_port, A2 
                           => n17081, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n84);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U7 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n58, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n52);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U5 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n56, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n51);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U10 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n53, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n48);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U6 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n2, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n46);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U40 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n115, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n5, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n59, C2 => 
                           n17297, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n116, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N119);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U41 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n8, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n31, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n10, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n81, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n12, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n80, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n116);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U56 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n20, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n5, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n21, C2 => 
                           n17297, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n22, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N112);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U57 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n8, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n23, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n10, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n24, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n12, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n25, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n22);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U48 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n4, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n5, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n6, C2 => 
                           n17297, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n7, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N114);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U49 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n8, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n9, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n10, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n11, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n12, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n13, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n7);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U50 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n64, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n5, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n71, C2 => 
                           n17737, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n148, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N115);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U51 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n8, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n30, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n10, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n31, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n12, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n81, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n148);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U60 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n14, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n5, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n15, C2 => 
                           n17297, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n16, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N113);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U61 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n8, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n17, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n10, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n18, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n12, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n19, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n16);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U70 : OAI21_X1 port map( B1 => n17112,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_C48_n110, A 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_n60, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N121);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U71 : OAI21_X1 port map( B1 => n17112,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_C48_n91, A 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_n60, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N122);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U64 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n32, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n40, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n91, C2 => 
                           n17737, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n92, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N106);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U65 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n12, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n9, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n43, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n93, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n10, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n35, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n92);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U172 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n46, B2 => 
                           n17077, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n48, C2 => 
                           n17102, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n98, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n93);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U173 : AOI22_X1 port map( A1 => n12649
                           , A2 => pipeline_stageE_EXE_ALU_alu_shift_C48_n51, 
                           B1 => pipeline_stageE_input1_to_ALU_1_port, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n52, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n98);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U96 : AOI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n13, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n73, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n11, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n1, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n108, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n91);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U98 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n105, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n72, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n84, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n74, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n109);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U76 : OAI21_X1 port map( B1 => n17112,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_C48_n27, A 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_n60, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N127);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U174 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n20, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n40, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n41, C2 => 
                           n17297, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n42, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N108);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U175 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n12, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n24, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n43, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n44, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n10, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n23, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n42);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U176 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n46, B2 => 
                           n17087, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n48, C2 => 
                           n17088, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n50, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n44);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U177 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_4_port, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n51, B1 => 
                           pipeline_stageE_input1_to_ALU_3_port, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n52, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n50);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U149 : OAI22_X1 port map( A1 => n17095
                           , A2 => pipeline_stageE_EXE_ALU_alu_shift_C48_n56, 
                           B1 => n17089, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n58, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n54);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U62 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n26, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n40, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n61, C2 => 
                           n17297, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n62, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N107);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U63 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n12, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n30, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n43, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n63, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n10, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n29, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n62);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U170 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n46, B2 => 
                           n17102, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n48, C2 => 
                           n17087, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n66, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n63);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U171 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_3_port, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n51, B1 => 
                           n12649, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n52, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n66);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U58 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n26, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n5, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n27, C2 => 
                           n17737, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n28, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N111);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U59 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n8, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n29, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n10, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n30, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n12, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n31, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n28);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U163 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_15_port, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n51, B1 => 
                           pipeline_stageE_input1_to_ALU_14_port, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n52, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n152);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U155 : OAI22_X1 port map( A1 => n17082
                           , A2 => pipeline_stageE_EXE_ALU_alu_shift_C48_n56, 
                           B1 => n17085, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n58, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n154);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U28 : AOI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n80, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n73, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n81, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n1, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n82, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n27);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U30 : AOI21_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n84, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n85, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n86, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n83);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U146 : OAI22_X1 port map( A1 => n17089
                           , A2 => pipeline_stageE_EXE_ALU_alu_shift_C48_n56, 
                           B1 => n17088, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n58, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n67);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U52 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n32, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n5, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n33, C2 => 
                           n17737, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n34, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N110);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U53 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n8, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n35, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n10, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n9, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n12, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n11, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n34);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U160 : OAI22_X1 port map( A1 => n17085
                           , A2 => pipeline_stageE_EXE_ALU_alu_shift_C48_n56, 
                           B1 => n17090, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n58, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n94);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U151 : OAI22_X1 port map( A1 => n17088
                           , A2 => pipeline_stageE_EXE_ALU_alu_shift_C48_n56, 
                           B1 => n17087, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n58, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n100);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U54 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n36, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n5, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n37, C2 => 
                           n17297, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n38, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N109);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U55 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n8, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n39, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n10, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n17, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n12, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n18, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n38);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U84 : OAI21_X1 port map( B1 => n17112,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_C48_n15, A 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_n60, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N129);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U34 : AOI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n76, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n73, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n77, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n1, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n75, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n15);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U43 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n111, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n40, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n112, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n5, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n113, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N120);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U46 : AOI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n12, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n78, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n10, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n79, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n114, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n113);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U38 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n99, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n5, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n68, C2 => 
                           n17737, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n118, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N118);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U39 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n8, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n11, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n10, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n13, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n12, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n74, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n118);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U137 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n46, B2 => 
                           n17097, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n48, C2 => 
                           n17118, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n127, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n11);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U138 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_18_port, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n51, B1 => 
                           pipeline_stageE_input1_to_ALU_17_port, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n52, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n127);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U166 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_14_port, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n51, B1 => 
                           pipeline_stageE_input1_to_ALU_13_port, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n52, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n133);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U72 : OAI21_X1 port map( B1 => n17112,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_C48_n61, A 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_n60, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N123);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U88 : AOI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n85, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n105, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n80, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n84, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n106, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n61);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U90 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n73, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n81, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n1, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n31, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n107);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U114 : OAI221_X1 port map( B1 => 
                           n17097, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n56, C1 => 
                           n17096, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n58, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n150, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n31);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U115 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_20_port, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n2, B1 => 
                           pipeline_stageE_input1_to_ALU_21_port, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n53, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n150);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U116 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n46, B2 => 
                           n17117, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n48, C2 => 
                           n17115, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n149, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n81);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U117 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_23_port, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n51, B1 => 
                           pipeline_stageE_input1_to_ALU_22_port, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n52, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n149);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U66 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n134, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n5, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n69, C2 => 
                           n17297, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n135, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N117);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U67 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n8, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n18, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n10, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n19, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n12, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n77, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n135);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U68 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n45, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n5, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n70, C2 => 
                           n17297, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n136, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N116);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U69 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n8, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n24, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n10, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n25, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n12, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n79, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n136);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U134 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n46, B2 => 
                           n17079, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n48, C2 => 
                           n17096, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n143, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n24);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U136 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_A_16_port, A2 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_n51, B1 => 
                           pipeline_stageE_input1_to_ALU_15_port, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n52, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n143);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U157 : OAI22_X1 port map( A1 => n17080
                           , A2 => pipeline_stageE_EXE_ALU_alu_shift_C48_n56, 
                           B1 => n17082, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n58, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n145);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U75 : OAI21_X1 port map( B1 => n17112,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_C48_n33, A 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_n60, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N126);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U25 : AOI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n74, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n73, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n13, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n1, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n87, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n33);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U27 : AOI21_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n84, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n72, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n86, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n88);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U131 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n46, B2 => 
                           n17092, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n48, C2 => 
                           n17117, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n124, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n13);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U133 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_22_port, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n51, B1 => 
                           pipeline_stageE_input1_to_ALU_21_port, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n52, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n124);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U74 : OAI21_X1 port map( B1 => n17112,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_C48_n37, A 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_n60, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N125);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U106 : AOI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n77, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n73, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n19, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n1, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n89, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n37);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U108 : AOI21_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n84, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n76, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n86, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n90);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U73 : OAI21_X1 port map( B1 => n17112,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_C48_n41, A 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_n60, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N124);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U103 : AOI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n79, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n73, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n25, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n1, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n101, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n41);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U105 : AOI21_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n84, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n78, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n86, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n102);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U42 : NOR2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n103, A2 => 
                           n17081, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n86);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U123 : OAI221_X1 port map( B1 => 
                           n17118, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n56, C1 => 
                           n17097, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n58, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n140, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n25);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U124 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_21_port, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n2, B1 => 
                           pipeline_stageE_input1_to_ALU_22_port, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n53, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n140);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U78 : OAI21_X1 port map( B1 => n17112,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_C48_n6, A =>
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n60, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N130);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U32 : AOI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n72, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n73, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n74, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n1, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n75, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n6);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U127 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n46, B2 => 
                           n17078, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n48, C2 => 
                           n17093, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n121, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n74);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U128 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_26_port, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n51, B1 => 
                           pipeline_stageE_input1_to_ALU_25_port, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n52, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n121);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U77 : OAI21_X1 port map( B1 => n17112,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_C48_n21, A 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_n60, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N128);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U31 : AOI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n78, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n73, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n79, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n1, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n75, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n21);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U125 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n46, B2 => 
                           n17115, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n48, C2 => 
                           n17086, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n139, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n79);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U126 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_24_port, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n51, B1 => 
                           pipeline_stageE_input1_to_ALU_23_port, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n52, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n139);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U79 : OAI21_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, B2 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_n71, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n60, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N131);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U33 : AOI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n85, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n73, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n80, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n1, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n75, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n71);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U143 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n46, B2 => 
                           n17093, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n48, C2 => 
                           n17094, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n153, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n80);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U144 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_27_port, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n51, B1 => 
                           pipeline_stageE_input1_to_ALU_26_port, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n52, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n153);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U80 : OAI21_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, B2 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_n70, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n60, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N132);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U35 : AOI21_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n78, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n1, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n117, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n70);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U141 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n46, B2 => 
                           n17094, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n48, C2 => 
                           n17083, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n144, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n78);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U142 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_28_port, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n51, B1 => 
                           pipeline_stageE_input1_to_ALU_27_port, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n52, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n144);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U83 : OAI21_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, B2 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_n69, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n60, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N133);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U37 : AOI21_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n76, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n1, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n117, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n69);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U81 : OAI21_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, B2 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_n68, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n60, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N134);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U17 : AOI21_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n72, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n1, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n117, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n68);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U24 : OAI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n58, A2 => 
                           n17094, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n56, B2 => 
                           n17083, C1 => n17303, C2 => n17104, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n72);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U82 : OAI21_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, B2 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_n59, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n60, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N135);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U3 : NAND2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, A2 
                           => pipeline_stageE_EXE_ALU_alu_shift_N136, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n60);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U36 : AOI21_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n85, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n1, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n117, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n59);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U109 : OAI21_X1 port map( B1 => n17081
                           , B2 => n17104, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n103, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n117);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U185 : NAND2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N136, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_3_port, ZN 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_n103);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U178 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n36, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n40, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n110, C2 => 
                           n17737, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n155, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N105);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U179 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n12, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n17, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n43, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n156, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n10, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n39, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n155);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U183 : OAI22_X1 port map( A1 => n17090
                           , A2 => pipeline_stageE_EXE_ALU_alu_shift_C48_n56, 
                           B1 => n17095, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n58, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n157);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U180 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n46, B2 => 
                           n17091, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n48, C2 => 
                           n17077, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n160, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n156);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U14 : NAND2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n1, A2 => 
                           n17302, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n5);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U169 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_13_port, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n51, B1 => 
                           pipeline_stageE_input1_to_ALU_12_port, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n52, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n162);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U99 : AOI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n19, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n73, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n18, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n1, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n163, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n110);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U101 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n105, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n76, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n84, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n77, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n164);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U129 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n46, B2 => 
                           n17086, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n48, C2 => 
                           n17078, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n165, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n77);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U130 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_25_port, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n51, B1 => 
                           pipeline_stageE_input1_to_ALU_24_port, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n52, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n165);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U118 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n46, B2 => 
                           n17083, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n48, C2 => 
                           n17104, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n166, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n76);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U119 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_29_port, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n51, B1 => 
                           pipeline_stageE_input1_to_ALU_28_port, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n52, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n166);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U139 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n46, B2 => 
                           n17096, C1 => n17097, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n48, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n167, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n18);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U140 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_17_port, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n51, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_A_16_port, B2 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_n52, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n167);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U120 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n56, B2 => 
                           n17084, C1 => n17118, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n58, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n169, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n19);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U122 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_22_port, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n2, B1 => 
                           pipeline_stageE_input1_to_ALU_23_port, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n53, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n169);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U18 : NAND2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n73, A2 => 
                           n17302, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n40);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U2 : NOR2_X1 port map( A1 => n17081, 
                           A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_3_port, ZN 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_n73);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U153 : OAI22_X1 port map( A1 => n17087
                           , A2 => pipeline_stageE_EXE_ALU_alu_shift_C48_n56, 
                           B1 => n17102, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n58, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n170);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U16 : NAND2_X1 port map( A1 => n17742,
                           A2 => n17303, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n58);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U9 : NAND2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, A2 
                           => n17303, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n56);
   pipeline_stageE_EXE_ALU_alu_shift_C48_U148 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_30_port, B => 
                           pipeline_stageE_EXE_ALU_alu_shift_N136, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n58, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n85);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U114 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n4, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n130);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U76 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n48, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n128);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U77 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n81, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n127);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U47 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n40, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n121);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U62 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n33, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n95);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U50 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n31, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n117);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U59 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n42, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n102);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U56 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n50, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n107);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U53 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n16, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n113);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U105 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n73, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n72);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U113 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n104, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n84);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U65 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n20, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n88);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U97 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n169, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n168);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U5 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n12, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n56);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U108 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n162, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n161);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U36 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n154, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n153);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U187 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n85, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n45);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U40 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n144, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n143);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U184 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n77, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n37);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U33 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n140, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n139);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U176 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n170, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n98);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U178 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n64, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n28);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U6 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n53, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n17);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U99 : AND2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_3_port, A2 
                           => n17302, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n131);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U101 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n135, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n134);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U112 : AND2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_3_port, A2 
                           => n17081, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n74);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U181 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n58, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n11);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U94 : OAI21_X1 port map( B1 => n17112,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_C86_n29, A 
                           => pipeline_stageE_EXE_ALU_alu_shift_C86_n4, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N216);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U87 : OAI21_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, B2 
                           => pipeline_stageE_EXE_ALU_alu_shift_C86_n6, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n4, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N209);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U82 : OAI21_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, B2 
                           => pipeline_stageE_EXE_ALU_alu_shift_C86_n3, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n4, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N211);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U84 : OAI21_X1 port map( B1 => n17112,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_C86_n61, A 
                           => pipeline_stageE_EXE_ALU_alu_shift_C86_n4, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N212);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U95 : OAI21_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, B2 
                           => pipeline_stageE_EXE_ALU_alu_shift_C86_n5, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n4, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N210);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U75 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n127, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n12, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n128, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n53, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n129, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N218);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U78 : AOI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n15, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n82, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n19, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n83, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n130, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n129);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U46 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n121, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n53, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n112, C2 => 
                           n17302, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n122, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N219);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U48 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n56, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n68, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n19, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n71, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n15, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n69, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n122);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U91 : OAI21_X1 port map( B1 => n17112,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_C86_n112, A 
                           => pipeline_stageE_EXE_ALU_alu_shift_C86_n4, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N203);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U42 : AOI21_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n75, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n1, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n109, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n112);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U61 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n95, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n53, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n7, C2 => 
                           n17302, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n96, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N224);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U63 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n56, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n31, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n19, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n63, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n15, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n97, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n96);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U90 : OAI21_X1 port map( B1 => n17112,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_C86_n10, A 
                           => pipeline_stageE_EXE_ALU_alu_shift_C86_n4, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N205);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U89 : OAI21_X1 port map( B1 => n17112,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_C86_n36, A 
                           => pipeline_stageE_EXE_ALU_alu_shift_C86_n4, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N204);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U88 : OAI21_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, B2 
                           => pipeline_stageE_EXE_ALU_alu_shift_C86_n7, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n4, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N208);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U30 : AOI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n98, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n70, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n99, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n1, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n84, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n7);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U85 : OAI21_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, B2 
                           => pipeline_stageE_EXE_ALU_alu_shift_C86_n8, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n4, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N207);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U86 : OAI21_X1 port map( B1 => n17112,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_C86_n9, A =>
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n4, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N206);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U73 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n45, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n53, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n5, C2 => 
                           n17302, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n80, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N226);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U74 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n56, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n50, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n19, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n48, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n15, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n81, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n80);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U38 : AOI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n82, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n70, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n83, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n1, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n84, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n5);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U93 : OAI21_X1 port map( B1 => n17112,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_C86_n13, A 
                           => pipeline_stageE_EXE_ALU_alu_shift_C86_n4, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N217);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U92 : OAI21_X1 port map( B1 => n17112,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_C86_n38, A 
                           => pipeline_stageE_EXE_ALU_alu_shift_C86_n4, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N215);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U49 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n117, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n53, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n36, C2 => 
                           n17302, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n118, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N220);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U51 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n56, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n63, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n19, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n97, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n15, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n99, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n118);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U43 : AOI21_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n98, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n1, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n109, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n36);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U81 : OAI21_X1 port map( B1 => n17112,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_C86_n46, A 
                           => pipeline_stageE_EXE_ALU_alu_shift_C86_n4, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N214);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U83 : OAI21_X1 port map( B1 => n17112,
                           B2 => pipeline_stageE_EXE_ALU_alu_shift_C86_n54, A 
                           => pipeline_stageE_EXE_ALU_alu_shift_C86_n4, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N213);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U58 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n102, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n53, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n8, C2 => 
                           n17302, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n103, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N223);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U60 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n56, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n40, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n19, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n68, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n15, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n71, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n103);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U29 : AOI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n75, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n70, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n69, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n1, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n84, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n8);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U55 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n107, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n53, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n9, C2 => 
                           n17302, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n108, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N222);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U57 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n56, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n48, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n19, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n81, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n15, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n83, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n108);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U45 : AOI21_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n82, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n1, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n109, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n9);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U52 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n113, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n53, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n10, C2 => 
                           n17302, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n114, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N221);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U54 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n56, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n57, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n19, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n90, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n15, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n92, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n114);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U44 : AOI21_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n91, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n1, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n109, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n10);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U110 : OAI21_X1 port map( B1 => n17119
                           , B2 => n17081, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n104, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n109);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U67 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n37, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n53, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n3, C2 => 
                           n17302, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n67, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N227);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U68 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n56, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n42, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n19, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n40, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n15, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n68, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n67);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U104 : AOI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n69, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n70, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n71, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n1, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n72, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n3);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U106 : AOI21_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n74, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n75, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n76, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n73);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U64 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n88, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n53, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n6, C2 => 
                           n17302, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n89, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N225);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U66 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n56, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n16, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n19, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n57, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n15, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n90, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n89);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U31 : AOI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n91, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n70, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n92, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n1, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n84, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n6);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U69 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n28, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n53, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n61, C2 => 
                           n17302, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n62, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N228);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U70 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n56, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n33, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n19, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n31, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n15, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n63, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n62);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U96 : AOI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n99, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n70, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n97, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n1, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n168, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n61);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U98 : AOI21_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n74, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n98, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n76, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n169);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U71 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n11, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n53, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n54, C2 => 
                           n17302, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n55, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N229);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U72 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n56, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n20, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n19, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n16, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n15, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n57, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n55);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U107 : AOI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n92, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n70, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n90, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n1, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n161, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n54);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U109 : AOI21_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n74, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n91, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n76, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n162);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U169 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n45, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n12, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n46, C2 => 
                           n17302, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n47, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N230);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U170 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n15, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n48, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n17, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n49, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n19, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n50, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n47);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U154 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n21, B2 => 
                           n17096, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n23, C2 => 
                           n17079, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n111, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n50);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U155 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_19_port, A2 => n17110,
                           B1 => pipeline_stageE_input1_to_ALU_20_port, B2 => 
                           n17111, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n111);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U171 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n21, B2 => 
                           n17086, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n23, C2 => 
                           n17115, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n52, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n49);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U172 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_27_port, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n26, B1 => 
                           pipeline_stageE_input1_to_ALU_28_port, B2 => n17111,
                           ZN => pipeline_stageE_EXE_ALU_alu_shift_C86_n52);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U138 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n21, B2 => 
                           n17100, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n23, C2 => 
                           n15425, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n133, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n48);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U139 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_15_port, A2 => n17110,
                           B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_A_16_port, B2 
                           => n17111, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n133);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U35 : AOI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n83, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n70, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n81, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n1, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n153, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n46);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U37 : AOI21_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n74, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n82, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n76, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n154);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U111 : NOR2_X1 port map( A1 => n17081,
                           A2 => pipeline_stageE_EXE_ALU_alu_shift_C86_n104, ZN
                           => pipeline_stageE_EXE_ALU_alu_shift_C86_n76);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U144 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n21, B2 => 
                           n17091, C1 => n17103, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n23, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n156, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n82);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U145 : AOI22_X1 port map( A1 => n17110
                           , A2 => pipeline_stageE_input1_to_ALU_3_port, B1 => 
                           pipeline_stageE_input1_to_ALU_4_port, B2 => n17111, 
                           ZN => pipeline_stageE_EXE_ALU_alu_shift_C86_n156);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U126 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n21, B2 => 
                           n17085, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n23, C2 => 
                           n17090, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n158, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n81);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U127 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_11_port, A2 => n17110,
                           B1 => pipeline_stageE_input1_to_ALU_12_port, B2 => 
                           n17111, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n158);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U120 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n21, B2 => 
                           n17088, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n23, C2 => 
                           n17087, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n160, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n83);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U121 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_7_port, A2 => n17110, 
                           B1 => pipeline_stageE_input1_to_ALU_8_port, B2 => 
                           n17111, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n160);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U188 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n21, B2 => 
                           n17116, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n23, C2 => 
                           n17084, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n87, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n85);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U189 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_23_port, A2 => n17110,
                           B1 => n17158, B2 => n17111, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n87);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U156 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n37, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n12, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n38, C2 => 
                           n17302, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n39, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N231);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U157 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n15, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n40, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n17, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n41, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n19, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n42, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n39);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U148 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n21, B2 => 
                           n17097, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n23, C2 => 
                           n17096, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n106, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n42);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U149 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_20_port, A2 => n17110,
                           B1 => pipeline_stageE_input1_to_ALU_21_port, B2 => 
                           n17111, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n106);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U158 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n21, B2 => 
                           n17078, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n23, C2 => 
                           n17086, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n44, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n41);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U159 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_28_port, A2 => n17110,
                           B1 => pipeline_stageE_input1_to_ALU_29_port, B2 => 
                           n17111, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n44);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U132 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n21, B2 => 
                           n17101, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n23, C2 => 
                           n17100, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n126, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n40);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U133 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_A_16_port, A2 
                           => n17110, B1 => 
                           pipeline_stageE_input1_to_ALU_17_port, B2 => n17111,
                           ZN => pipeline_stageE_EXE_ALU_alu_shift_C86_n126);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U39 : AOI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n75, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n136, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n69, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n74, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n143, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n38);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U41 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n70, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n71, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n1, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n68, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n144);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U174 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n21, B2 => 
                           n17082, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n23, C2 => 
                           n17085, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n146, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n68);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U175 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_12_port, A2 => n17110,
                           B1 => pipeline_stageE_input1_to_ALU_13_port, B2 => 
                           n17111, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n146);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U116 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n21, B2 => 
                           n17089, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n23, C2 => 
                           n17088, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n149, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n71);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U117 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_8_port, A2 => n17110, 
                           B1 => pipeline_stageE_input1_to_ALU_9_port, B2 => 
                           n17111, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n149);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U146 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n21, B2 => 
                           n17077, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n23, C2 => 
                           n17091, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n152, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n69);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U147 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_4_port, A2 => n17110, 
                           B1 => pipeline_stageE_input1_to_ALU_5_port, B2 => 
                           n17111, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n152);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U185 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n21, B2 => 
                           n17092, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n23, C2 => 
                           n17116, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n79, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n77);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U186 : AOI22_X1 port map( A1 => n17158
                           , A2 => n17110, B1 => n17159, B2 => n17111, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n79);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U160 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n28, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n12, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n29, C2 => 
                           n17302, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n30, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N232);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U161 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n15, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n31, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n17, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n32, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n19, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n33, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n30);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U150 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n21, B2 => 
                           n17118, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n23, C2 => 
                           n17097, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n101, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n33);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U151 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_21_port, A2 => n17110,
                           B1 => pipeline_stageE_input1_to_ALU_22_port, B2 => 
                           n17111, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n101);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U162 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n21, B2 => 
                           n17093, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n23, C2 => 
                           n17078, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n35, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n32);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U163 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_29_port, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n26, B1 => 
                           pipeline_stageE_input1_to_ALU_30_port, B2 => n17111,
                           ZN => pipeline_stageE_EXE_ALU_alu_shift_C86_n35);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U134 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n21, B2 => 
                           n17738, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n23, C2 => 
                           n17101, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n120, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n31);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U135 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_17_port, A2 => n17110,
                           B1 => pipeline_stageE_input1_to_ALU_18_port, B2 => 
                           n17111, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n120);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U32 : AOI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n97, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n70, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n63, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n1, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n139, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n29);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U34 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n136, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n98, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n74, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n99, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n140);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U122 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n21, B2 => 
                           n17102, C1 => n17077, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n23, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n172, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n99);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U123 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_5_port, A2 => n17110, 
                           B1 => pipeline_stageE_input1_to_ALU_6_port, B2 => 
                           n17111, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n172);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U140 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n21, B2 => 
                           n17080, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n23, C2 => 
                           n17082, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n142, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n63);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U141 : AOI22_X1 port map( A1 => n17160
                           , A2 => n17110, B1 => 
                           pipeline_stageE_input1_to_ALU_14_port, B2 => n17111,
                           ZN => pipeline_stageE_EXE_ALU_alu_shift_C86_n142);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U128 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n21, B2 => 
                           n17095, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n23, C2 => 
                           n17089, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n171, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n97);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U129 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_9_port, A2 => n17110, 
                           B1 => pipeline_stageE_input1_to_ALU_10_port, B2 => 
                           n17111, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n171);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U179 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n21, B2 => 
                           n17117, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n23, C2 => 
                           n17092, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n66, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n64);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U180 : AOI22_X1 port map( A1 => n17159
                           , A2 => n17110, B1 => 
                           pipeline_stageE_input1_to_ALU_26_port, B2 => n17111,
                           ZN => pipeline_stageE_EXE_ALU_alu_shift_C86_n66);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U164 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n11, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n12, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n13, C2 => 
                           n17302, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n14, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N233);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U166 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n15, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n16, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n17, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n18, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n19, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n20, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n14);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U152 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n21, B2 => 
                           n17084, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n23, C2 => 
                           n17118, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n94, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n20);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U153 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_22_port, A2 => n17110,
                           B1 => pipeline_stageE_input1_to_ALU_23_port, B2 => 
                           n17111, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n94);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U167 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n21, B2 => 
                           n17094, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n23, C2 => 
                           n17093, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n25, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n18);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U173 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_30_port, A2 => n17110,
                           B1 => pipeline_stageE_EXE_ALU_alu_shift_N136, B2 => 
                           n17111, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n25);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U14 : NAND2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n1, A2 => 
                           n17302, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n53);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U136 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n21, B2 => 
                           n17079, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n23, C2 => 
                           n17738, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n116, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n16);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U137 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_18_port, A2 => n17110,
                           B1 => pipeline_stageE_input1_to_ALU_19_port, B2 => 
                           n17111, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n116);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U100 : AOI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n90, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n70, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n57, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n1, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n134, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n13);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U102 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n136, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n91, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n74, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n92, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n135);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U124 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n21, B2 => 
                           n17087, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n23, C2 => 
                           n17102, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n167, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n92);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U125 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_6_port, A2 => n17110, 
                           B1 => pipeline_stageE_input1_to_ALU_7_port, B2 => 
                           n17111, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n167);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U118 : OAI221_X1 port map( B1 => 
                           n17103, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n21, C1 => 
                           n17119, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n23, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n163, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n91);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U119 : AOI22_X1 port map( A1 => n17110
                           , A2 => n12649, B1 => 
                           pipeline_stageE_input1_to_ALU_3_port, B2 => n17111, 
                           ZN => pipeline_stageE_EXE_ALU_alu_shift_C86_n163);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U142 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n21, B2 => 
                           n15425, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n23, C2 => 
                           n17080, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n138, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n57);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U143 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_14_port, A2 => n17110,
                           B1 => pipeline_stageE_input1_to_ALU_15_port, B2 => 
                           n17111, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n138);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U130 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n21, B2 => 
                           n17090, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n23, C2 => 
                           n17095, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n165, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n90);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U131 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_10_port, A2 => n17110,
                           B1 => pipeline_stageE_input1_to_ALU_11_port, B2 => 
                           n17111, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n165);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U15 : NAND2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n70, A2 => 
                           n17302, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n12);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U2 : NOR2_X1 port map( A1 => n17081, 
                           A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_3_port, ZN 
                           => pipeline_stageE_EXE_ALU_alu_shift_C86_n70);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U182 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n21, B2 => 
                           n17115, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n23, C2 => 
                           n17117, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n60, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n58);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U183 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_26_port, A2 => n17110,
                           B1 => pipeline_stageE_input1_to_ALU_27_port, B2 => 
                           n17111, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n60);
   pipeline_stageE_EXE_ALU_alu_shift_C86_U165 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_N202, B => 
                           pipeline_stageE_input1_to_ALU_1_port, S => n17111, Z
                           => pipeline_stageE_EXE_ALU_alu_shift_C86_n75);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M0_0_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_N202, B => 
                           pipeline_stageE_EXE_ALU_alu_shift_N136, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_0_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_0_1 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_1_port, B => 
                           pipeline_stageE_EXE_ALU_alu_shift_N202, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_1_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_0_2 : MUX2_X1 port map( A => n12649
                           , B => pipeline_stageE_input1_to_ALU_1_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_2_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_0_3 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_3_port, B => n12649, S
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, 
                           Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_3_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_0_5 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_5_port, B => 
                           pipeline_stageE_input1_to_ALU_4_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_5_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_0_6 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_6_port, B => 
                           pipeline_stageE_input1_to_ALU_5_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_6_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_0_7 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_7_port, B => 
                           pipeline_stageE_input1_to_ALU_6_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_7_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_0_8 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_8_port, B => 
                           pipeline_stageE_input1_to_ALU_7_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_8_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_0_9 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_9_port, B => 
                           pipeline_stageE_input1_to_ALU_8_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_9_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_0_10 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_10_port, B => 
                           pipeline_stageE_input1_to_ALU_9_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_10_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_0_11 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_11_port, B => 
                           pipeline_stageE_input1_to_ALU_10_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_11_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_0_12 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_12_port, B => 
                           pipeline_stageE_input1_to_ALU_11_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_12_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_0_13 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_13_port, B => 
                           pipeline_stageE_input1_to_ALU_12_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_13_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_0_14 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_14_port, B => 
                           pipeline_stageE_input1_to_ALU_13_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_14_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_0_15 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_15_port, B => 
                           pipeline_stageE_input1_to_ALU_14_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_15_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_0_16 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_A_16_port, B 
                           => pipeline_stageE_input1_to_ALU_15_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_16_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_0_17 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_17_port, B => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_A_16_port, S 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, 
                           Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_17_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_0_18 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_18_port, B => 
                           pipeline_stageE_input1_to_ALU_17_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_18_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_0_19 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_19_port, B => 
                           pipeline_stageE_input1_to_ALU_18_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_19_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_0_20 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_20_port, B => 
                           pipeline_stageE_input1_to_ALU_19_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_20_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_0_21 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_21_port, B => 
                           pipeline_stageE_input1_to_ALU_20_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_21_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_0_22 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_22_port, B => 
                           pipeline_stageE_input1_to_ALU_21_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_22_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_0_23 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_23_port, B => 
                           pipeline_stageE_input1_to_ALU_22_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_23_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_0_24 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_24_port, B => 
                           pipeline_stageE_input1_to_ALU_23_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_24_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_0_25 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_25_port, B => 
                           pipeline_stageE_input1_to_ALU_24_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_25_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_0_26 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_26_port, B => 
                           pipeline_stageE_input1_to_ALU_25_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_26_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_0_27 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_27_port, B => 
                           pipeline_stageE_input1_to_ALU_26_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_27_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_0_28 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_28_port, B => 
                           pipeline_stageE_input1_to_ALU_27_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_28_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_0_29 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_29_port, B => 
                           pipeline_stageE_input1_to_ALU_28_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_29_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_0_30 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_30_port, B => 
                           pipeline_stageE_input1_to_ALU_29_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_30_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_0_31 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_N136, B => 
                           pipeline_stageE_input1_to_ALU_30_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_31_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M0_1_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_0_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_30_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_0_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M0_1_1 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_1_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_31_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_1_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_1_2 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_2_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_0_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_2_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_1_3 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_3_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_1_port, S 
                           => n17298, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_3_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_1_4 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_4_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_2_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_4_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_1_5 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_5_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_3_port, S 
                           => n17298, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_5_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_1_6 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_6_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_4_port, S 
                           => n17298, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_6_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_1_7 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_7_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_5_port, S 
                           => n17298, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_7_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_1_8 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_8_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_6_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_8_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_1_9 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_9_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_7_port, S 
                           => n17298, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_9_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_1_10 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_10_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_8_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_10_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_1_11 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_11_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_9_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_11_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_1_12 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_12_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_10_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_12_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_1_13 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_13_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_11_port, S 
                           => n17298, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_13_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_1_14 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_14_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_12_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_14_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_1_15 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_15_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_13_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_15_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_1_16 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_16_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_14_port, S 
                           => n17298, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_16_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_1_17 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_17_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_15_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_17_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_1_18 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_18_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_16_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_18_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_1_19 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_19_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_17_port, S 
                           => n17298, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_19_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_1_20 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_20_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_18_port, S 
                           => n17298, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_20_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_1_21 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_21_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_19_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_21_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_1_22 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_22_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_20_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_22_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_1_23 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_23_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_21_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_23_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_1_24 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_24_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_22_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_24_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_1_25 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_25_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_23_port, S 
                           => n17298, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_25_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_1_26 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_26_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_24_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_26_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_1_27 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_27_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_25_port, S 
                           => n17298, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_27_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_1_28 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_28_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_26_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_28_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_1_29 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_29_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_27_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_29_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_1_30 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_30_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_28_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_30_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_1_31 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_31_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_1_29_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_31_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M0_2_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_0_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_28_port, S 
                           => n17114, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_0_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M0_2_1 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_1_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_29_port, S 
                           => n17114, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_1_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M0_2_2 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_2_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_30_port, S 
                           => n17114, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_2_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M0_2_3 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_3_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_31_port, S 
                           => n17114, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_3_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_2_4 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_4_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_0_port, S 
                           => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_4_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_2_5 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_5_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_1_port, S 
                           => n17114, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_5_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_2_6 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_6_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_2_port, S 
                           => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_6_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_2_7 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_7_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_3_port, S 
                           => n17114, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_7_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_2_8 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_8_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_4_port, S 
                           => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_8_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_2_9 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_9_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_5_port, S 
                           => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_9_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_2_10 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_10_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_6_port, S 
                           => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_10_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_2_11 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_11_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_7_port, S 
                           => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_11_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_2_12 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_12_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_8_port, S 
                           => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_12_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_2_13 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_13_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_9_port, S 
                           => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_13_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_2_14 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_14_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_10_port, S 
                           => n17114, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_14_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_2_15 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_15_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_11_port, S 
                           => n17114, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_15_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_2_16 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_16_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_12_port, S 
                           => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_16_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_2_17 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_17_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_13_port, S 
                           => n17114, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_17_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_2_18 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_18_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_14_port, S 
                           => n17114, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_18_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_2_19 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_19_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_15_port, S 
                           => n17114, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_19_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_2_20 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_20_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_16_port, S 
                           => n17114, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_20_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_2_21 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_21_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_17_port, S 
                           => n17114, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_21_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_2_22 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_22_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_18_port, S 
                           => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_22_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_2_23 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_23_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_19_port, S 
                           => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_23_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_2_24 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_24_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_20_port, S 
                           => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_24_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_2_25 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_25_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_21_port, S 
                           => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_25_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_2_26 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_26_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_22_port, S 
                           => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_26_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_2_27 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_27_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_23_port, S 
                           => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_27_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_2_28 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_28_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_24_port, S 
                           => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_28_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_2_29 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_29_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_25_port, S 
                           => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_29_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_2_30 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_30_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_26_port, S 
                           => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_30_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_2_31 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_31_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_2_27_port, S 
                           => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_31_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M0_3_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_0_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_24_port, S 
                           => n17301, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_0_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M0_3_1 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_1_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_25_port, S 
                           => n17301, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_1_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M0_3_2 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_2_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_26_port, S 
                           => n17301, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_2_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M0_3_3 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_3_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_27_port, S 
                           => n17301, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_3_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M0_3_4 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_4_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_28_port, S 
                           => n17301, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_4_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M0_3_5 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_5_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_29_port, S 
                           => n17301, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_5_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M0_3_6 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_6_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_30_port, S 
                           => n17301, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_6_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M0_3_7 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_7_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_31_port, S 
                           => n17301, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_7_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_3_8 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_8_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_0_port, S 
                           => n17301, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_8_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_3_9 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_9_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_1_port, S 
                           => n17301, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_9_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_3_10 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_10_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_2_port, S 
                           => n17301, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_10_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_3_11 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_11_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_3_port, S 
                           => n17301, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_11_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_3_12 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_12_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_4_port, S 
                           => n17300, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_12_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_3_13 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_13_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_5_port, S 
                           => n17300, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_13_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_3_14 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_14_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_6_port, S 
                           => n17300, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_14_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_3_15 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_15_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_7_port, S 
                           => n17300, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_15_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_3_16 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_16_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_8_port, S 
                           => n17300, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_16_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_3_17 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_17_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_9_port, S 
                           => n17300, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_17_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_3_18 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_18_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_10_port, S 
                           => n17300, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_18_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_3_19 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_19_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_11_port, S 
                           => n17300, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_19_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_3_20 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_20_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_12_port, S 
                           => n17300, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_20_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_3_21 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_21_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_13_port, S 
                           => n17300, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_21_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_3_22 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_22_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_14_port, S 
                           => n17300, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_22_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_3_23 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_23_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_15_port, S 
                           => n17300, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_23_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_3_24 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_24_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_16_port, S 
                           => n17301, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_24_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_3_25 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_25_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_17_port, S 
                           => n17300, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_25_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_3_26 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_26_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_18_port, S 
                           => n17300, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_26_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_3_27 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_27_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_19_port, S 
                           => n17299, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_27_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_3_28 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_28_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_20_port, S 
                           => n17299, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_28_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_3_29 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_29_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_21_port, S 
                           => n17299, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_29_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_3_30 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_30_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_22_port, S 
                           => n17299, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_30_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_3_31 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_31_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_3_23_port, S 
                           => n17300, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_31_port);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M0_4_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_0_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_16_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N39);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M0_4_1 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_1_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_17_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N40);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M0_4_2 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_2_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_18_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N41);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M0_4_3 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_3_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_19_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N42);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M0_4_4 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_4_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_20_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N43);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M0_4_5 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_5_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_21_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N44);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M0_4_6 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_6_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_22_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N45);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M0_4_7 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_7_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_23_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N46);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M0_4_8 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_8_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_24_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N47);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M0_4_9 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_9_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_25_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N48);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M0_4_10 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_10_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_26_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N49);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M0_4_11 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_11_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_27_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N50);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M0_4_12 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_12_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_28_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N51);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M0_4_13 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_13_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_29_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N52);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M0_4_14 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_14_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_30_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N53);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M0_4_15 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_15_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_31_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N54);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_4_16 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_16_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_0_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N55);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_4_17 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_17_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_1_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N56);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_4_18 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_18_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_2_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N57);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_4_19 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_19_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_3_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N58);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_4_20 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_20_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_4_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N59);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_4_21 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_21_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_5_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N60);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_4_22 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_22_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_6_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N61);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_4_23 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_23_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_7_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N62);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_4_24 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_24_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_8_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N63);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_4_25 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_25_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_9_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N64);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_4_26 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_26_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_10_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N65);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_4_27 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_27_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_11_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N66);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_4_28 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_28_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_12_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N67);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_4_29 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_29_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_13_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N68);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_4_30 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_30_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_14_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N69);
   pipeline_stageE_EXE_ALU_alu_shift_C10_M1_4_31 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_31_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C10_ML_int_4_15_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N70);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_0_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_N202, B => 
                           pipeline_stageE_input1_to_ALU_1_port, S => n17113, Z
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_0_port
                           );
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_0_1_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_1_port, B => n12649, S
                           => n17113, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_1_port
                           );
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_0_2_0 : MUX2_X1 port map( A => 
                           n12649, B => pipeline_stageE_input1_to_ALU_3_port, S
                           => n17113, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_2_port
                           );
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_0_3_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_3_port, B => 
                           pipeline_stageE_input1_to_ALU_4_port, S => n17113, Z
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_3_port
                           );
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_0_4_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_4_port, B => 
                           pipeline_stageE_input1_to_ALU_5_port, S => n17113, Z
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_4_port
                           );
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_0_5_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_5_port, B => 
                           pipeline_stageE_input1_to_ALU_6_port, S => n17113, Z
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_5_port
                           );
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_0_6_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_6_port, B => 
                           pipeline_stageE_input1_to_ALU_7_port, S => n17113, Z
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_6_port
                           );
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_0_7_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_7_port, B => 
                           pipeline_stageE_input1_to_ALU_8_port, S => n17113, Z
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_7_port
                           );
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_0_8_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_8_port, B => 
                           pipeline_stageE_input1_to_ALU_9_port, S => n17113, Z
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_8_port
                           );
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_0_9_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_9_port, B => 
                           pipeline_stageE_input1_to_ALU_10_port, S => n17113, 
                           Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_9_port
                           );
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_0_10_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_10_port, B => 
                           pipeline_stageE_input1_to_ALU_11_port, S => n17113, 
                           Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_10_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_0_11_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_11_port, B => 
                           pipeline_stageE_input1_to_ALU_12_port, S => n17113, 
                           Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_11_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_0_12_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_12_port, B => 
                           pipeline_stageE_input1_to_ALU_13_port, S => n17113, 
                           Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_12_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_0_13_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_13_port, B => 
                           pipeline_stageE_input1_to_ALU_14_port, S => n17113, 
                           Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_13_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_0_14_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_14_port, B => 
                           pipeline_stageE_input1_to_ALU_15_port, S => n17113, 
                           Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_14_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_0_15_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_15_port, B => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_A_16_port, S 
                           => n17113, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_15_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_0_16_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_A_16_port, B 
                           => pipeline_stageE_input1_to_ALU_17_port, S => 
                           n17113, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_16_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_0_17_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_17_port, B => 
                           pipeline_stageE_input1_to_ALU_18_port, S => n17113, 
                           Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_17_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_0_18_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_18_port, B => 
                           pipeline_stageE_input1_to_ALU_19_port, S => n17113, 
                           Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_18_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_0_19_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_19_port, B => 
                           pipeline_stageE_input1_to_ALU_20_port, S => n17113, 
                           Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_19_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_0_20_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_20_port, B => 
                           pipeline_stageE_input1_to_ALU_21_port, S => n17113, 
                           Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_20_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_0_21_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_21_port, B => 
                           pipeline_stageE_input1_to_ALU_22_port, S => n17113, 
                           Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_21_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_0_22_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_22_port, B => 
                           pipeline_stageE_input1_to_ALU_23_port, S => n17113, 
                           Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_22_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_0_23_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_23_port, B => 
                           pipeline_stageE_input1_to_ALU_24_port, S => n17113, 
                           Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_23_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_0_24_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_24_port, B => 
                           pipeline_stageE_input1_to_ALU_25_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_24_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_0_25_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_25_port, B => 
                           pipeline_stageE_input1_to_ALU_26_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_25_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_0_26_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_26_port, B => 
                           pipeline_stageE_input1_to_ALU_27_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_26_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_0_27_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_27_port, B => 
                           pipeline_stageE_input1_to_ALU_28_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_27_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_0_28_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_28_port, B => 
                           pipeline_stageE_input1_to_ALU_29_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_28_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_0_29_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_29_port, B => 
                           pipeline_stageE_input1_to_ALU_30_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_29_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_0_30_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_30_port, B => 
                           pipeline_stageE_EXE_ALU_alu_shift_N136, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_30_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_0_31_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_N136, B => 
                           pipeline_stageE_EXE_ALU_alu_shift_N202, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_31_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_1_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_0_port
                           , B => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_2_port
                           , S => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_0_port
                           );
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_1_1 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_1_port
                           , B => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_3_port
                           , S => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_1_port
                           );
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_1_2_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_2_port
                           , B => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_4_port
                           , S => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_2_port
                           );
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_1_3_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_3_port
                           , B => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_5_port
                           , S => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_3_port
                           );
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_1_4_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_4_port
                           , B => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_6_port
                           , S => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_4_port
                           );
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_1_5_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_5_port
                           , B => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_7_port
                           , S => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_5_port
                           );
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_1_6_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_6_port
                           , B => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_8_port
                           , S => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_6_port
                           );
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_1_7_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_7_port
                           , B => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_9_port
                           , S => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_7_port
                           );
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_1_8_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_8_port
                           , B => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_10_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_8_port
                           );
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_1_9_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_9_port
                           , B => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_11_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_9_port
                           );
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_1_10_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_10_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_12_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_10_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_1_11_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_11_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_13_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_11_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_1_12_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_12_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_14_port, S 
                           => n17298, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_12_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_1_13_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_13_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_15_port, S 
                           => n17298, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_13_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_1_14_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_14_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_16_port, S 
                           => n17298, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_14_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_1_15_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_15_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_17_port, S 
                           => n17298, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_15_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_1_16_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_16_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_18_port, S 
                           => n17298, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_16_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_1_17_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_17_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_19_port, S 
                           => n17298, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_17_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_1_18_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_18_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_20_port, S 
                           => n17298, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_18_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_1_19_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_19_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_21_port, S 
                           => n17298, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_19_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_1_20_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_20_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_22_port, S 
                           => n17298, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_20_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_1_21_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_21_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_23_port, S 
                           => n17298, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_21_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_1_22_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_22_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_24_port, S 
                           => n17298, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_22_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_1_23_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_23_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_25_port, S 
                           => n17298, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_23_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_1_24_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_24_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_26_port, S 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_SH_1_port, 
                           Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_24_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_1_25_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_25_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_27_port, S 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_SH_1_port, 
                           Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_25_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_1_26_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_26_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_28_port, S 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_SH_1_port, 
                           Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_26_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_1_27_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_27_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_29_port, S 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_SH_1_port, 
                           Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_27_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_1_28_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_28_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_30_port, S 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_SH_1_port, 
                           Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_28_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_1_29_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_29_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_31_port, S 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_SH_1_port, 
                           Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_29_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_1_30_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_30_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_0_port
                           , S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_1_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_30_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_1_31_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_31_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_1_1_port
                           , S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_1_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_31_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_2_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_0_port
                           , B => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_4_port
                           , S => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_0_port
                           );
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_2_1 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_1_port
                           , B => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_5_port
                           , S => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_1_port
                           );
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_2_2 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_2_port
                           , B => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_6_port
                           , S => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_2_port
                           );
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_2_3 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_3_port
                           , B => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_7_port
                           , S => n17114, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_3_port
                           );
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_2_4_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_4_port
                           , B => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_8_port
                           , S => n17114, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_4_port
                           );
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_2_5_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_5_port
                           , B => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_9_port
                           , S => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_5_port
                           );
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_2_6_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_6_port
                           , B => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_10_port, S 
                           => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_6_port
                           );
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_2_7_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_7_port
                           , B => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_11_port, S 
                           => n17114, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_7_port
                           );
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_2_8_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_8_port
                           , B => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_12_port, S 
                           => n17114, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_8_port
                           );
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_2_9_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_9_port
                           , B => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_13_port, S 
                           => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_9_port
                           );
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_2_10_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_10_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_14_port, S 
                           => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_10_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_2_11_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_11_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_15_port, S 
                           => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_11_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_2_12_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_12_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_16_port, S 
                           => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_12_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_2_13_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_13_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_17_port, S 
                           => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_13_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_2_14_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_14_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_18_port, S 
                           => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_14_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_2_15_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_15_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_19_port, S 
                           => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_15_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_2_16_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_16_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_20_port, S 
                           => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_16_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_2_17_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_17_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_21_port, S 
                           => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_17_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_2_18_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_18_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_22_port, S 
                           => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_18_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_2_19_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_19_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_23_port, S 
                           => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_19_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_2_20_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_20_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_24_port, S 
                           => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_20_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_2_21_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_21_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_25_port, S 
                           => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_21_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_2_22_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_22_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_26_port, S 
                           => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_22_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_2_23_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_23_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_27_port, S 
                           => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_23_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_2_24_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_24_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_28_port, S 
                           => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_24_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_2_25_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_25_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_29_port, S 
                           => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_25_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_2_26_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_26_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_30_port, S 
                           => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_26_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_2_27_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_27_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_31_port, S 
                           => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_27_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_2_28_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_28_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_0_port
                           , S => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_28_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_2_29_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_29_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_1_port
                           , S => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_29_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_2_30_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_30_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_2_port
                           , S => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_30_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_2_31_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_31_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_2_3_port
                           , S => n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_31_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_3_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_0_port
                           , B => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_8_port
                           , S => n17299, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_0_port
                           );
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_3_1 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_1_port
                           , B => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_9_port
                           , S => n17299, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_1_port
                           );
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_3_2 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_2_port
                           , B => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_10_port, S 
                           => n17299, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_2_port
                           );
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_3_3 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_3_port
                           , B => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_11_port, S 
                           => n17299, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_3_port
                           );
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_3_4 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_4_port
                           , B => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_12_port, S 
                           => n17299, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_4_port
                           );
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_3_5 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_5_port
                           , B => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_13_port, S 
                           => n17299, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_5_port
                           );
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_3_6 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_6_port
                           , B => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_14_port, S 
                           => n17299, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_6_port
                           );
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_3_7 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_7_port
                           , B => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_15_port, S 
                           => n17299, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_7_port
                           );
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_3_8_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_8_port
                           , B => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_16_port, S 
                           => n17299, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_8_port
                           );
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_3_9_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_9_port
                           , B => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_17_port, S 
                           => n17299, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_9_port
                           );
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_3_10_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_10_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_18_port, S 
                           => n17299, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_10_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_3_11_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_11_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_19_port, S 
                           => n17299, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_11_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_3_12_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_12_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_20_port, S 
                           => n17296, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_12_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_3_13_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_13_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_21_port, S 
                           => n17296, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_13_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_3_14_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_14_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_22_port, S 
                           => n17296, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_14_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_3_15_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_15_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_23_port, S 
                           => n17296, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_15_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_3_16_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_16_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_24_port, S 
                           => n17296, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_16_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_3_17_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_17_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_25_port, S 
                           => n17296, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_17_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_3_18_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_18_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_26_port, S 
                           => n17296, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_18_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_3_19_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_19_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_27_port, S 
                           => n17296, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_19_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_3_20_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_20_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_28_port, S 
                           => n17296, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_20_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_3_21_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_21_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_29_port, S 
                           => n17296, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_21_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_3_22_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_22_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_30_port, S 
                           => n17296, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_22_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_3_23_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_23_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_31_port, S 
                           => n17296, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_23_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_3_24_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_24_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_0_port
                           , S => n17300, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_24_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_3_25_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_25_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_1_port
                           , S => n17299, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_25_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_3_26_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_26_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_2_port
                           , S => n17301, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_26_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_3_27_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_27_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_3_port
                           , S => n17301, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_27_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_3_28_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_28_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_4_port
                           , S => n17296, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_28_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_3_29_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_29_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_5_port
                           , S => n17296, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_29_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_3_30_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_30_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_6_port
                           , S => n17301, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_30_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_3_31_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_31_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_3_7_port
                           , S => n17299, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_31_port);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_4_0 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_0_port
                           , B => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_16_port, S 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, 
                           Z => pipeline_stageE_EXE_ALU_alu_shift_N7);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_4_1 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_1_port
                           , B => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_17_port, S 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, 
                           Z => pipeline_stageE_EXE_ALU_alu_shift_N8);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_4_2 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_2_port
                           , B => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_18_port, S 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, 
                           Z => pipeline_stageE_EXE_ALU_alu_shift_N9);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_4_3 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_3_port
                           , B => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_19_port, S 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, 
                           Z => pipeline_stageE_EXE_ALU_alu_shift_N10);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_4_4 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_4_port
                           , B => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_20_port, S 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, 
                           Z => pipeline_stageE_EXE_ALU_alu_shift_N11);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_4_5 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_5_port
                           , B => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_21_port, S 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, 
                           Z => pipeline_stageE_EXE_ALU_alu_shift_N12);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_4_6 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_6_port
                           , B => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_22_port, S 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, 
                           Z => pipeline_stageE_EXE_ALU_alu_shift_N13);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_4_7 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_7_port
                           , B => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_23_port, S 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, 
                           Z => pipeline_stageE_EXE_ALU_alu_shift_N14);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_4_8 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_8_port
                           , B => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_24_port, S 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, 
                           Z => pipeline_stageE_EXE_ALU_alu_shift_N15);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_4_9 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_9_port
                           , B => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_25_port, S 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, 
                           Z => pipeline_stageE_EXE_ALU_alu_shift_N16);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_4_10 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_10_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_26_port, S 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, 
                           Z => pipeline_stageE_EXE_ALU_alu_shift_N17);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_4_11 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_11_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_27_port, S 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, 
                           Z => pipeline_stageE_EXE_ALU_alu_shift_N18);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_4_12 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_12_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_28_port, S 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, 
                           Z => pipeline_stageE_EXE_ALU_alu_shift_N19);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_4_13 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_13_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_29_port, S 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, 
                           Z => pipeline_stageE_EXE_ALU_alu_shift_N20);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_4_14 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_14_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_30_port, S 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, 
                           Z => pipeline_stageE_EXE_ALU_alu_shift_N21);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_4_15 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_15_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_31_port, S 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, 
                           Z => pipeline_stageE_EXE_ALU_alu_shift_N22);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_4_16 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_16_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_0_port
                           , S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, Z 
                           => pipeline_stageE_EXE_ALU_alu_shift_N23);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_4_17 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_17_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_1_port
                           , S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, Z 
                           => pipeline_stageE_EXE_ALU_alu_shift_N24);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_4_18 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_18_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_2_port
                           , S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, Z 
                           => pipeline_stageE_EXE_ALU_alu_shift_N25);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_4_19 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_19_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_3_port
                           , S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, Z 
                           => pipeline_stageE_EXE_ALU_alu_shift_N26);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_4_20 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_20_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_4_port
                           , S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, Z 
                           => pipeline_stageE_EXE_ALU_alu_shift_N27);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_4_21 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_21_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_5_port
                           , S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, Z 
                           => pipeline_stageE_EXE_ALU_alu_shift_N28);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_4_22 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_22_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_6_port
                           , S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, Z 
                           => pipeline_stageE_EXE_ALU_alu_shift_N29);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_4_23 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_23_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_7_port
                           , S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, Z 
                           => pipeline_stageE_EXE_ALU_alu_shift_N30);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_4_24 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_24_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_8_port
                           , S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, Z 
                           => pipeline_stageE_EXE_ALU_alu_shift_N31);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_4_25 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_25_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_9_port
                           , S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, Z 
                           => pipeline_stageE_EXE_ALU_alu_shift_N32);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_4_26 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_26_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_10_port, S 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, 
                           Z => pipeline_stageE_EXE_ALU_alu_shift_N33);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_4_27 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_27_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_11_port, S 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, 
                           Z => pipeline_stageE_EXE_ALU_alu_shift_N34);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_4_28 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_28_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_12_port, S 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, 
                           Z => pipeline_stageE_EXE_ALU_alu_shift_N35);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_4_29 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_29_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_13_port, S 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, 
                           Z => pipeline_stageE_EXE_ALU_alu_shift_N36);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_4_30 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_30_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_14_port, S 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, 
                           Z => pipeline_stageE_EXE_ALU_alu_shift_N37);
   pipeline_stageE_EXE_ALU_alu_shift_C8_M1_4_31 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_31_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C8_MR_int_4_15_port, S 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, 
                           Z => pipeline_stageE_EXE_ALU_alu_shift_N38);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U87 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n28, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n101);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U88 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n29, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n100);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U107 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n94, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n93);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U100 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n43, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n21);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U96 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n63, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n27);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U97 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n2, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n33);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U84 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n23, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n96);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U80 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n7, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n104);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U81 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n9, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n103);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U110 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n91, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n90);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U101 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n121, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N149);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U104 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n123, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n122);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U8 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n38, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n6);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U99 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n22, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n97);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U44 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n89, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n69);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U112 : AND2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n68, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n41, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N165);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U46 : AND2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n67, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n41, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N166);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U47 : AND2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n59, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n41, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N167);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U48 : AND2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n41, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n58, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N168);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U98 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n12, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n37);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U5 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n3, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n41);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U59 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n156, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n155);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U9 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n50, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n57);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U7 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n49, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n55);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U11 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n44, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n51);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U86 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n100, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n38, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n101, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n3, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n102, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N151);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U89 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n10, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n78, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n99, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n59, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n8, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n79, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n102);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U70 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n18, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n3, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n19, C2 => 
                           n17297, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n20, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N144);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U71 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n6, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n21, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n8, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n22, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n10, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n23, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n20);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U62 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n2, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n3, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n4, C2 => 
                           n17297, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n5, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N146);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U63 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n6, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n7, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n8, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n9, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n10, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n11, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n5);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U64 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n63, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n3, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n70, C2 => 
                           n17297, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n138, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N147);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U65 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n6, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n28, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n8, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n29, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n10, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n79, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n138);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U74 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n12, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n3, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n13, C2 => 
                           n17297, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n14, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N145);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U75 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n6, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n15, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n8, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n16, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n10, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n17, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n14);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U37 : NOR2_X1 port map( A1 => n17112, 
                           A2 => pipeline_stageE_EXE_ALU_alu_shift_C50_n95, ZN 
                           => pipeline_stageE_EXE_ALU_alu_shift_N153);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U38 : NOR2_X1 port map( A1 => n17112, 
                           A2 => pipeline_stageE_EXE_ALU_alu_shift_C50_n80, ZN 
                           => pipeline_stageE_EXE_ALU_alu_shift_N154);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U166 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n30, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n38, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n80, C2 => 
                           n17297, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n81, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N138);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U167 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n10, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n7, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n41, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n82, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n8, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n33, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n81);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U168 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n44, B2 => 
                           n17102, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n21, C2 => 
                           n17077, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n87, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n82);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U169 : AOI22_X1 port map( A1 => n12649
                           , A2 => pipeline_stageE_EXE_ALU_alu_shift_C86_n26, 
                           B1 => pipeline_stageE_input1_to_ALU_1_port, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n27, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n87);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U106 : AOI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n11, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n73, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n9, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n72, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n93, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n80);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U108 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n92, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n67, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n76, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n71, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n94);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U33 : NOR2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, A2 
                           => pipeline_stageE_EXE_ALU_alu_shift_C50_n25, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N159);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U162 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n18, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n38, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n39, C2 => 
                           n17297, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n40, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N140);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U163 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n10, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n22, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n41, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n42, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n8, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n21, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n40);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U164 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n44, B2 => 
                           n17088, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n21, C2 => 
                           n17087, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n48, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n42);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U165 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_4_port, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n26, B1 => 
                           pipeline_stageE_input1_to_ALU_3_port, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n27, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n48);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U178 : AOI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n51, B2 => 
                           pipeline_stageE_input1_to_ALU_10_port, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n167, C2 => 
                           pipeline_stageE_input1_to_ALU_9_port, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n53, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n18);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U179 : OAI22_X1 port map( A1 => n17095
                           , A2 => pipeline_stageE_EXE_ALU_alu_shift_C50_n55, 
                           B1 => n17089, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n57, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n53);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U158 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n24, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n38, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n60, C2 => 
                           n17297, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n61, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N139);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U159 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n10, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n28, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n41, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n62, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n8, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n27, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n61);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U160 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n44, B2 => 
                           n17087, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n21, C2 => 
                           n17102, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n65, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n62);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U161 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_3_port, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n26, B1 => 
                           n12649, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n50, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n65);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U72 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n24, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n3, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n25, C2 => 
                           n17297, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n26, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N143);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U73 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n6, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n27, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n8, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n28, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n10, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n29, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n26);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U127 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n44, B2 => 
                           n17079, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n21, C2 => 
                           n17738, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n142, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n28);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U128 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_15_port, A2 => n17110,
                           B1 => pipeline_stageE_input1_to_ALU_14_port, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n50, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n142);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U148 : OAI22_X1 port map( A1 => n17082
                           , A2 => pipeline_stageE_EXE_ALU_alu_shift_C50_n55, 
                           B1 => n17085, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n57, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n144);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U55 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n78, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n73, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n59, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n76, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n79, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n72, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n25);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U176 : AOI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n51, B2 => 
                           pipeline_stageE_input1_to_ALU_9_port, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n167, C2 => 
                           pipeline_stageE_input1_to_ALU_8_port, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n66, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n24);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U177 : OAI22_X1 port map( A1 => n17089
                           , A2 => pipeline_stageE_EXE_ALU_alu_shift_C50_n55, 
                           B1 => n17088, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n57, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n66);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U66 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n30, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n3, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n31, C2 => 
                           n17297, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n32, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N142);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U67 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n6, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n33, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n8, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n7, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n10, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n9, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n32);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U149 : AOI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n51, B2 => 
                           pipeline_stageE_input1_to_ALU_12_port, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n167, C2 => 
                           pipeline_stageE_input1_to_ALU_11_port, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n83, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n2);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U150 : OAI22_X1 port map( A1 => n17085
                           , A2 => pipeline_stageE_EXE_ALU_alu_shift_C50_n55, 
                           B1 => n17090, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n57, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n83);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U180 : AOI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n51, B2 => 
                           pipeline_stageE_input1_to_ALU_8_port, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n167, C2 => 
                           pipeline_stageE_input1_to_ALU_7_port, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n88, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n30);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U181 : OAI22_X1 port map( A1 => n17088
                           , A2 => pipeline_stageE_EXE_ALU_alu_shift_C50_n55, 
                           B1 => n17087, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n57, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n88);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U68 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n34, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n3, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n35, C2 => 
                           n17297, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n36, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N141);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U69 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n6, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n37, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n8, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n15, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n10, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n16, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n36);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U40 : NOR2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, A2 
                           => pipeline_stageE_EXE_ALU_alu_shift_C50_n13, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N161);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U92 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n74, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n72, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n68, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n73, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n13);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U83 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n96, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n38, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n97, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n3, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n98, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N152);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U85 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n10, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n75, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n99, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n58, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n8, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n77, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n98);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U79 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n103, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n38, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n104, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n3, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n105, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N150);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U82 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n10, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n71, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n99, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n67, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n8, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n11, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n105);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U125 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n44, B2 => 
                           n17738, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n46, C2 => 
                           n17101, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n117, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n7);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U126 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_14_port, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n26, B1 => 
                           n17160, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n50, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n117);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U119 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n44, B2 => 
                           n17118, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n21, C2 => 
                           n17097, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n120, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n9);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U120 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_18_port, A2 => n17110,
                           B1 => pipeline_stageE_input1_to_ALU_17_port, B2 => 
                           n17111, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n120);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U39 : NOR2_X1 port map( A1 => n17112, 
                           A2 => pipeline_stageE_EXE_ALU_alu_shift_C50_n60, ZN 
                           => pipeline_stageE_EXE_ALU_alu_shift_N155);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U109 : AOI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n79, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n73, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n29, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n72, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n90, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n60);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U111 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n92, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n59, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n76, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n78, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n91);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U121 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n44, B2 => 
                           n17084, C1 => n17118, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n46, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n141, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n29);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U122 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n49, A2 => 
                           pipeline_stageE_input1_to_ALU_19_port, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n50, B2 => 
                           pipeline_stageE_input1_to_ALU_18_port, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n141);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U141 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n44, B2 => 
                           n17115, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n21, C2 => 
                           n17117, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n139, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n79);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U142 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_23_port, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n49, B1 => 
                           pipeline_stageE_input1_to_ALU_22_port, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n50, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n139);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U103 : AOI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n16, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n6, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n15, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n41, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n122, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n121);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U105 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n10, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n74, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n99, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n68, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n8, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n17, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n123);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U13 : NOR2_X1 port map( A1 => n17297, 
                           A2 => pipeline_stageE_EXE_ALU_alu_shift_C50_n124, ZN
                           => pipeline_stageE_EXE_ALU_alu_shift_C50_n99);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U76 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n97, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n38, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n43, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n3, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n125, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N148);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U77 : AOI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n10, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n77, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n8, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n23, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n126, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n125);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U78 : NOR3_X1 port map( A1 => n17297, 
                           A2 => n17296, A3 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n69, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n126);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U154 : OAI22_X1 port map( A1 => n17080
                           , A2 => pipeline_stageE_EXE_ALU_alu_shift_C50_n55, 
                           B1 => n17082, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n57, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n132);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U151 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n44, B2 => 
                           n17096, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n21, C2 => 
                           n17079, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n137, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n22);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U152 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_A_16_port, A2 
                           => n17110, B1 => 
                           pipeline_stageE_input1_to_ALU_15_port, B2 => n17111,
                           ZN => pipeline_stageE_EXE_ALU_alu_shift_C50_n137);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U32 : NOR2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, A2 
                           => pipeline_stageE_EXE_ALU_alu_shift_C50_n31, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N158);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U54 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n71, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n73, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n67, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n76, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n11, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n72, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n31);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U138 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n44, B2 => 
                           n17117, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n46, C2 => 
                           n17092, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n108, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n11);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U140 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_22_port, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n49, B1 => 
                           pipeline_stageE_input1_to_ALU_21_port, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n50, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n108);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U31 : NOR2_X1 port map( A1 => n17112, 
                           A2 => pipeline_stageE_EXE_ALU_alu_shift_C50_n35, ZN 
                           => pipeline_stageE_EXE_ALU_alu_shift_N157);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U53 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n74, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n73, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n68, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n76, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n17, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n72, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n35);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U36 : NOR2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, A2 
                           => pipeline_stageE_EXE_ALU_alu_shift_C50_n39, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N156);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U57 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n23, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n72, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n77, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n73, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n89, C2 => 
                           n17296, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n39);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U117 : OAI221_X1 port map( B1 => 
                           n17118, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n55, C1 => 
                           n17097, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n57, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n128, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n23);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U118 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_22_port, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n51, B1 => 
                           pipeline_stageE_input1_to_ALU_21_port, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n167, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n128);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U35 : NOR2_X1 port map( A1 => n17112, 
                           A2 => pipeline_stageE_EXE_ALU_alu_shift_C50_n4, ZN 
                           => pipeline_stageE_EXE_ALU_alu_shift_N162);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U90 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n71, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n72, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n67, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n73, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n4);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U132 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n44, B2 => 
                           n17093, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n46, C2 => 
                           n17078, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n114, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n71);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U133 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_26_port, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n49, B1 => 
                           pipeline_stageE_input1_to_ALU_25_port, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n50, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n114);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U34 : NOR2_X1 port map( A1 => n17112, 
                           A2 => pipeline_stageE_EXE_ALU_alu_shift_C50_n19, ZN 
                           => pipeline_stageE_EXE_ALU_alu_shift_N160);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U56 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n75, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n73, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n58, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n76, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n77, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n72, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n19);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U145 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n44, B2 => 
                           n17086, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n46, C2 => 
                           n17115, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n131, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n77);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U146 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_24_port, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n49, B1 => 
                           pipeline_stageE_input1_to_ALU_23_port, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n50, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n131);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U41 : NOR2_X1 port map( A1 => n17112, 
                           A2 => pipeline_stageE_EXE_ALU_alu_shift_C50_n70, ZN 
                           => pipeline_stageE_EXE_ALU_alu_shift_N163);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U91 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n78, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n72, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n59, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n73, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n70);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U134 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n44, B2 => 
                           n17094, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n46, C2 => 
                           n17093, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n143, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n78);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U135 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_27_port, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n49, B1 => 
                           pipeline_stageE_input1_to_ALU_26_port, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n50, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n143);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U15 : NOR3_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n69, A2 => 
                           n17112, A3 => n17296, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N164);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U156 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n44, B2 => 
                           n17083, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n21, C2 => 
                           n17094, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n127, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n75);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U157 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_28_port, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n49, B1 => 
                           pipeline_stageE_input1_to_ALU_27_port, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n27, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n127);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U51 : OAI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n55, A2 => 
                           n17083, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n46, B2 => 
                           n17104, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n57, C2 => 
                           n17094, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n67);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U52 : OAI22_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n57, A2 => 
                           n17083, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n55, B2 => 
                           n17104, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n59);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U93 : NOR2_X1 port map( A1 => n17104, 
                           A2 => pipeline_stageE_EXE_ALU_alu_shift_C50_n57, ZN 
                           => pipeline_stageE_EXE_ALU_alu_shift_C50_n58);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U170 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n34, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n38, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n95, C2 => 
                           n17297, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n145, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N137);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U171 : AOI222_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n10, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n15, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n41, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n146, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n8, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n37, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n145);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U174 : AOI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n51, B2 => 
                           pipeline_stageE_input1_to_ALU_11_port, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n167, C2 => 
                           pipeline_stageE_input1_to_ALU_10_port, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n147, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n12);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U175 : OAI22_X1 port map( A1 => n17090
                           , A2 => pipeline_stageE_EXE_ALU_alu_shift_C50_n55, 
                           B1 => n17095, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n57, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n147);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U172 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n44, B2 => 
                           n17077, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n46, C2 => 
                           n17091, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n151, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n146);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U6 : NAND2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n72, A2 => 
                           n17297, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n3);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U129 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n44, B2 => 
                           n17101, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n46, C2 => 
                           n17100, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n153, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n15);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U131 : AOI22_X1 port map( A1 => n17160
                           , A2 => pipeline_stageE_EXE_ALU_alu_shift_C50_n49, 
                           B1 => pipeline_stageE_input1_to_ALU_12_port, B2 => 
                           n17111, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n153);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U28 : NOR2_X1 port map( A1 => n17739, 
                           A2 => n17112, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n148);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U58 : AOI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n17, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n73, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n16, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n72, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n155, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n95);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U60 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n92, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n68, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n76, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n74, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n156);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U136 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n44, B2 => 
                           n17078, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n46, C2 => 
                           n17086, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n157, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n74);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U137 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_25_port, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n49, B1 => 
                           pipeline_stageE_input1_to_ALU_24_port, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n50, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n157);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U115 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n44, B2 => 
                           n17104, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n21, C2 => 
                           n17083, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n158, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n68);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U116 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_29_port, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n49, B1 => 
                           pipeline_stageE_input1_to_ALU_28_port, B2 => n17111,
                           ZN => pipeline_stageE_EXE_ALU_alu_shift_C50_n158);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U23 : NOR2_X1 port map( A1 => n17081, 
                           A2 => n17739, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n92);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U27 : NAND2_X1 port map( A1 => n17081,
                           A2 => n17739, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n124);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U123 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n44, B2 => 
                           n17097, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n21, C2 => 
                           n17096, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n159, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n16);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U124 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_17_port, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n49, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_A_16_port, B2 
                           => pipeline_stageE_EXE_ALU_alu_shift_C50_n50, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n159);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U143 : OAI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n55, B2 => 
                           n17084, C1 => n17118, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n57, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n160, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n17);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U144 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_input1_to_ALU_23_port, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n51, B1 => 
                           pipeline_stageE_input1_to_ALU_22_port, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n167, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n160);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U12 : NAND2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n73, A2 => 
                           n17297, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n38);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U182 : AOI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n51, B2 => 
                           pipeline_stageE_input1_to_ALU_7_port, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n167, C2 => 
                           pipeline_stageE_input1_to_ALU_6_port, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n161, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n34);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U183 : OAI22_X1 port map( A1 => n17087
                           , A2 => pipeline_stageE_EXE_ALU_alu_shift_C50_n55, 
                           B1 => n17102, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n57, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n161);
   pipeline_stageE_EXE_ALU_alu_shift_C50_U102 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n75, B => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n58, S => 
                           n17074, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n89);
   pipeline_stageE_EXE_ALU_alu_shift_C88_U38 : AND2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_14_port, 
                           A2 => n17737, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N248);
   pipeline_stageE_EXE_ALU_alu_shift_C88_U33 : AND2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_9_port, 
                           A2 => n17297, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N243);
   pipeline_stageE_EXE_ALU_alu_shift_C88_U35 : AND2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_10_port, 
                           A2 => n17302, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N244);
   pipeline_stageE_EXE_ALU_alu_shift_C88_U39 : AND2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_8_port, 
                           A2 => n17302, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N242);
   pipeline_stageE_EXE_ALU_alu_shift_C88_U13 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_n10, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_0_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_U10 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_n9, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_1_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_U16 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_n4, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_6_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_U37 : AND2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_15_port, 
                           A2 => n17302, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N249);
   pipeline_stageE_EXE_ALU_alu_shift_C88_U36 : AND2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_13_port, 
                           A2 => n17297, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N247);
   pipeline_stageE_EXE_ALU_alu_shift_C88_U11 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_n8, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_2_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_U32 : AND2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_12_port, 
                           A2 => n17302, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N246);
   pipeline_stageE_EXE_ALU_alu_shift_C88_U34 : AND2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_11_port, 
                           A2 => n17297, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N245);
   pipeline_stageE_EXE_ALU_alu_shift_C88_U15 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_n5, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_5_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_U14 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_n6, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_4_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_U12 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_n7, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_3_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_U29 : AND2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_1_port, 
                           A2 => n17081, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_1_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_U17 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_n3, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_7_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_U30 : AND2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_2_port, 
                           A2 => n17081, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_2_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_U31 : AND2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_3_port, 
                           A2 => n17081, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_3_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_U46 : AND2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_1_port, 
                           A2 => n17303, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_1_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_U44 : AND2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_0_port, 
                           A2 => n17081, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_0_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_U48 : AND2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_0_port, 
                           A2 => n17303, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_0_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_U6 : NOR2_X1 port map( A1 => n17112, 
                           A2 => pipeline_stageE_EXE_ALU_alu_shift_C88_n3, ZN 
                           => pipeline_stageE_EXE_ALU_alu_shift_N241);
   pipeline_stageE_EXE_ALU_alu_shift_C88_U18 : NOR2_X1 port map( A1 => n17112, 
                           A2 => pipeline_stageE_EXE_ALU_alu_shift_C88_n9, ZN 
                           => pipeline_stageE_EXE_ALU_alu_shift_N235);
   pipeline_stageE_EXE_ALU_alu_shift_C88_U28 : NAND2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_1_port, 
                           A2 => n17739, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_n9);
   pipeline_stageE_EXE_ALU_alu_shift_C88_U9 : NOR2_X1 port map( A1 => n17112, 
                           A2 => pipeline_stageE_EXE_ALU_alu_shift_C88_n7, ZN 
                           => pipeline_stageE_EXE_ALU_alu_shift_N237);
   pipeline_stageE_EXE_ALU_alu_shift_C88_U8 : NOR2_X1 port map( A1 => n17112, 
                           A2 => pipeline_stageE_EXE_ALU_alu_shift_C88_n8, ZN 
                           => pipeline_stageE_EXE_ALU_alu_shift_N236);
   pipeline_stageE_EXE_ALU_alu_shift_C88_U7 : NOR2_X1 port map( A1 => n17112, 
                           A2 => pipeline_stageE_EXE_ALU_alu_shift_C88_n4, ZN 
                           => pipeline_stageE_EXE_ALU_alu_shift_N240);
   pipeline_stageE_EXE_ALU_alu_shift_C88_U25 : NAND2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_6_port, 
                           A2 => n17739, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_n4);
   pipeline_stageE_EXE_ALU_alu_shift_C88_U4 : NOR2_X1 port map( A1 => n17112, 
                           A2 => pipeline_stageE_EXE_ALU_alu_shift_C88_n5, ZN 
                           => pipeline_stageE_EXE_ALU_alu_shift_N239);
   pipeline_stageE_EXE_ALU_alu_shift_C88_U5 : NOR2_X1 port map( A1 => n17112, 
                           A2 => pipeline_stageE_EXE_ALU_alu_shift_C88_n6, ZN 
                           => pipeline_stageE_EXE_ALU_alu_shift_N238);
   pipeline_stageE_EXE_ALU_alu_shift_C88_U26 : NAND2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_2_port, 
                           A2 => n17739, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_n8);
   pipeline_stageE_EXE_ALU_alu_shift_C88_U22 : NAND2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_5_port, 
                           A2 => n17739, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_n5);
   pipeline_stageE_EXE_ALU_alu_shift_C88_U23 : NAND2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_4_port, 
                           A2 => n17739, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_n6);
   pipeline_stageE_EXE_ALU_alu_shift_C88_U27 : NAND2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_3_port, 
                           A2 => n17739, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_n7);
   pipeline_stageE_EXE_ALU_alu_shift_C88_U24 : NAND2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_7_port, 
                           A2 => n17739, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_n3);
   pipeline_stageE_EXE_ALU_alu_shift_C88_U19 : NOR2_X1 port map( A1 => n17112, 
                           A2 => pipeline_stageE_EXE_ALU_alu_shift_C88_n10, ZN 
                           => pipeline_stageE_EXE_ALU_alu_shift_N234);
   pipeline_stageE_EXE_ALU_alu_shift_C88_U43 : NAND2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_0_port, 
                           A2 => n17739, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_n10);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_0_1 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_1_port, B => 
                           pipeline_stageE_EXE_ALU_alu_shift_N202, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_1_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_0_2 : MUX2_X1 port map( A => n12649
                           , B => pipeline_stageE_input1_to_ALU_1_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_2_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_0_3 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_3_port, B => n12649, S
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, 
                           Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_3_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_0_4 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_4_port, B => 
                           pipeline_stageE_input1_to_ALU_3_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_4_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_0_5 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_5_port, B => 
                           pipeline_stageE_input1_to_ALU_4_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_5_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_0_6 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_6_port, B => 
                           pipeline_stageE_input1_to_ALU_5_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_6_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_0_7 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_7_port, B => 
                           pipeline_stageE_input1_to_ALU_6_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_7_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_0_8 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_8_port, B => 
                           pipeline_stageE_input1_to_ALU_7_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_8_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_0_9 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_9_port, B => 
                           pipeline_stageE_input1_to_ALU_8_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_9_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_0_10 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_10_port, B => 
                           pipeline_stageE_input1_to_ALU_9_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_10_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_0_11 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_11_port, B => 
                           pipeline_stageE_input1_to_ALU_10_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_11_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_0_12 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_12_port, B => 
                           pipeline_stageE_input1_to_ALU_11_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_12_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_0_13 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_13_port, B => 
                           pipeline_stageE_input1_to_ALU_12_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_13_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_0_14 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_14_port, B => 
                           pipeline_stageE_input1_to_ALU_13_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_14_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_0_15 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_15_port, B => 
                           pipeline_stageE_input1_to_ALU_14_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_15_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_0_16 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_A_16_port, B 
                           => pipeline_stageE_input1_to_ALU_15_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_16_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_0_17 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_17_port, B => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_A_16_port, S 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, 
                           Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_17_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_0_18 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_18_port, B => 
                           pipeline_stageE_input1_to_ALU_17_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_18_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_0_19 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_19_port, B => 
                           pipeline_stageE_input1_to_ALU_18_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_19_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_0_20 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_20_port, B => 
                           pipeline_stageE_input1_to_ALU_19_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_20_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_0_21 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_21_port, B => 
                           pipeline_stageE_input1_to_ALU_20_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_21_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_0_22 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_22_port, B => 
                           pipeline_stageE_input1_to_ALU_21_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_22_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_0_23 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_23_port, B => 
                           pipeline_stageE_input1_to_ALU_22_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_23_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_0_24 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_24_port, B => 
                           pipeline_stageE_input1_to_ALU_23_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_24_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_0_25 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_25_port, B => 
                           pipeline_stageE_input1_to_ALU_24_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_25_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_0_26 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_26_port, B => 
                           pipeline_stageE_input1_to_ALU_25_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_26_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_0_27 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_27_port, B => 
                           pipeline_stageE_input1_to_ALU_26_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_27_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_0_28 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_28_port, B => 
                           pipeline_stageE_input1_to_ALU_27_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_28_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_0_29 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_29_port, B => 
                           pipeline_stageE_input1_to_ALU_28_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_29_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_0_30 : MUX2_X1 port map( A => 
                           pipeline_stageE_input1_to_ALU_30_port, B => 
                           pipeline_stageE_input1_to_ALU_29_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_30_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_0_31 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_N136, B => 
                           pipeline_stageE_input1_to_ALU_30_port, S => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_31_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_1_2 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_2_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_0_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_2_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_1_3 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_3_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_1_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_3_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_1_4 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_4_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_2_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_4_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_1_5 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_5_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_3_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_5_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_1_6 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_6_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_4_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_6_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_1_7 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_7_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_5_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_7_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_1_8 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_8_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_6_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_8_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_1_9 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_9_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_7_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_9_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_1_10 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_10_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_8_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_10_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_1_11 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_11_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_9_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_11_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_1_12 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_12_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_10_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_12_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_1_13 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_13_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_11_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_13_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_1_14 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_14_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_12_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_14_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_1_15 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_15_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_13_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_15_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_1_16 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_16_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_14_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_16_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_1_17 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_17_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_15_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_17_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_1_18 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_18_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_16_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_18_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_1_19 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_19_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_17_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_19_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_1_20 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_20_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_18_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_20_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_1_21 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_21_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_19_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_21_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_1_22 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_22_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_20_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_22_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_1_23 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_23_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_21_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_23_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_1_24 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_24_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_22_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_24_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_1_25 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_25_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_23_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_25_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_1_26 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_26_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_24_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_26_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_1_27 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_27_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_25_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_27_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_1_28 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_28_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_26_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_28_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_1_29 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_29_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_27_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_29_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_1_30 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_30_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_28_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_30_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_1_31 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_31_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_29_port, S 
                           => n17099, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_31_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_2_4 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_4_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_0_port, S 
                           => n17114, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_4_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_2_5 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_5_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_1_port, S 
                           => n17114, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_5_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_2_6 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_6_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_2_port, S 
                           => n17114, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_6_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_2_7 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_7_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_3_port, S 
                           => n17114, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_7_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_2_8 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_8_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_4_port, S 
                           => n17114, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_8_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_2_9 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_9_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_5_port, S 
                           => n17114, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_9_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_2_10 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_10_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_6_port, S 
                           => n17114, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_10_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_2_11 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_11_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_7_port, S 
                           => n17114, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_11_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_2_12 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_12_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_8_port, S 
                           => n17114, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_12_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_2_13 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_13_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_9_port, S 
                           => n17114, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_13_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_2_14 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_14_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_10_port, S 
                           => n17114, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_14_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_2_15 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_15_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_11_port, S 
                           => n17114, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_15_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_2_16 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_16_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_12_port, S 
                           => n17114, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_16_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_2_17 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_17_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_13_port, S 
                           => n17114, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_17_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_2_18 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_18_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_14_port, S 
                           => n17114, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_18_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_2_19 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_19_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_15_port, S 
                           => n17114, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_19_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_2_20 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_20_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_16_port, S 
                           => n17114, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_20_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_2_21 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_21_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_17_port, S 
                           => n17114, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_21_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_2_22 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_22_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_18_port, S 
                           => n17114, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_22_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_2_23 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_23_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_19_port, S 
                           => n17114, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_23_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_2_24 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_24_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_20_port, S 
                           => n17114, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_24_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_2_25 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_25_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_21_port, S 
                           => n17114, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_25_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_2_26 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_26_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_22_port, S 
                           => n17114, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_26_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_2_27 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_27_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_23_port, S 
                           => n17114, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_27_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_2_28 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_28_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_24_port, S 
                           => n17114, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_28_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_2_29 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_29_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_25_port, S 
                           => n17114, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_29_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_2_30 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_30_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_26_port, S 
                           => n17114, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_30_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_2_31 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_31_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_2_27_port, S 
                           => n17114, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_31_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_3_8 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_8_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_0_port, S 
                           => n17296, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_8_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_3_9 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_9_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_1_port, S 
                           => n17301, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_9_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_3_10 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_10_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_2_port, S 
                           => n17300, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_10_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_3_11 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_11_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_3_port, S 
                           => n17301, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_11_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_3_12 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_12_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_4_port, S 
                           => n17301, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_12_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_3_13 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_13_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_5_port, S 
                           => n17300, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_13_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_3_14 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_14_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_6_port, S 
                           => n17300, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_14_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_3_15 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_15_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_7_port, S 
                           => n17299, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_15_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_3_16 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_16_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_8_port, S 
                           => n17296, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_16_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_3_17 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_17_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_9_port, S 
                           => n17299, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_17_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_3_18 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_18_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_10_port, S 
                           => n17301, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_18_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_3_19 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_19_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_11_port, S 
                           => n17296, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_19_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_3_20 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_20_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_12_port, S 
                           => n17300, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_20_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_3_21 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_21_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_13_port, S 
                           => n17296, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_21_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_3_22 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_22_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_14_port, S 
                           => n17300, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_22_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_3_23 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_23_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_15_port, S 
                           => n17301, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_23_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_3_24 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_24_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_16_port, S 
                           => n17301, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_24_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_3_25 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_25_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_17_port, S 
                           => n17299, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_25_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_3_26 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_26_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_18_port, S 
                           => n17300, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_26_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_3_27 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_27_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_19_port, S 
                           => n17296, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_27_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_3_28 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_28_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_20_port, S 
                           => n17300, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_28_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_3_29 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_29_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_21_port, S 
                           => n17301, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_29_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_3_30 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_30_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_22_port, S 
                           => n17299, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_30_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_3_31 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_31_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_3_23_port, S 
                           => n17299, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_31_port);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_4_16 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_16_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_0_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N250);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_4_17 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_17_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_1_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N251);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_4_18 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_18_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_2_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N252);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_4_19 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_19_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_3_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N253);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_4_20 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_20_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_4_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N254);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_4_21 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_21_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_5_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N255);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_4_22 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_22_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_6_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N256);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_4_23 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_23_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_7_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N257);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_4_24 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_24_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_8_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N258);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_4_25 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_25_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_9_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N259);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_4_26 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_26_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_10_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N260);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_4_27 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_27_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_11_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N261);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_4_28 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_28_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_12_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N262);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_4_29 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_29_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_13_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N263);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_4_30 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_30_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_14_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N264);
   pipeline_stageE_EXE_ALU_alu_shift_C88_M1_4_31 : MUX2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_31_port, B 
                           => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_4_15_port, S 
                           => n17112, Z => 
                           pipeline_stageE_EXE_ALU_alu_shift_N265);
   pipeline_stageD_evaluate_jump_target_add_29_U41 : INV_X1 port map( A => 
                           pipeline_stageD_offset_to_jump_temp_24_port, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n168);
   pipeline_stageD_evaluate_jump_target_add_29_U57 : INV_X1 port map( A => 
                           pipeline_stageD_offset_to_jump_temp_20_port, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n180);
   pipeline_stageD_evaluate_jump_target_add_29_U75 : INV_X1 port map( A => 
                           pipeline_stageD_offset_to_jump_temp_16_port, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n194);
   pipeline_stageD_evaluate_jump_target_add_29_U67 : INV_X1 port map( A => 
                           pipeline_stageD_offset_to_jump_temp_18_port, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n188);
   pipeline_stageD_evaluate_jump_target_add_29_U49 : INV_X1 port map( A => 
                           pipeline_stageD_offset_to_jump_temp_22_port, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n174);
   pipeline_stageD_evaluate_jump_target_add_29_U59 : XNOR2_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_add_29_n183, B 
                           => pipeline_stageD_evaluate_jump_target_add_29_n184,
                           ZN => pipeline_stageD_evaluate_jump_target_N34);
   pipeline_stageD_evaluate_jump_target_add_29_U14 : XNOR2_X1 port map( A => 
                           pipeline_nextPC_IFID_DEC_3_port, B => 
                           pipeline_stageD_offset_to_jump_temp_3_port, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n144);
   pipeline_stageD_evaluate_jump_target_add_29_U10 : XNOR2_X1 port map( A => 
                           pipeline_nextPC_IFID_DEC_5_port, B => 
                           pipeline_stageD_offset_to_jump_temp_5_port, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n138);
   pipeline_stageD_evaluate_jump_target_add_29_U12 : AOI22_X1 port map( A1 => 
                           pipeline_nextPC_IFID_DEC_4_port, A2 => 
                           pipeline_stageD_offset_to_jump_temp_4_port, B1 => 
                           n17412, B2 => n17455, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n141);
   pipeline_stageD_evaluate_jump_target_add_29_U8 : AOI22_X1 port map( A1 => 
                           pipeline_nextPC_IFID_DEC_6_port, A2 => 
                           pipeline_stageD_offset_to_jump_temp_6_port, B1 => 
                           n17361, B2 => n17456, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n135);
   pipeline_stageD_evaluate_jump_target_add_29_U6 : XNOR2_X1 port map( A => 
                           pipeline_nextPC_IFID_DEC_7_port, B => 
                           pipeline_stageD_offset_to_jump_temp_7_port, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n132);
   pipeline_stageD_evaluate_jump_target_add_29_U4 : AOI22_X1 port map( A1 => 
                           pipeline_nextPC_IFID_DEC_8_port, A2 => 
                           pipeline_stageD_offset_to_jump_temp_8_port, B1 => 
                           n17428, B2 => n17457, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n129);
   pipeline_stageD_evaluate_jump_target_add_29_U2 : XNOR2_X1 port map( A => 
                           pipeline_stageD_offset_to_jump_temp_9_port, B => 
                           pipeline_nextPC_IFID_DEC_9_port, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n126);
   pipeline_stageD_evaluate_jump_target_add_29_U97 : AOI22_X1 port map( A1 => 
                           pipeline_nextPC_IFID_DEC_10_port, A2 => 
                           pipeline_stageD_offset_to_jump_temp_10_port, B1 => 
                           n17440, B2 => n17458, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n213);
   pipeline_stageD_evaluate_jump_target_add_29_U93 : XNOR2_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_add_29_n209, B 
                           => n17174, ZN => 
                           pipeline_stageD_evaluate_jump_target_N44);
   pipeline_stageD_evaluate_jump_target_add_29_U95 : XNOR2_X1 port map( A => 
                           pipeline_nextPC_IFID_DEC_11_port, B => 
                           pipeline_stageD_offset_to_jump_temp_11_port, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n209);
   pipeline_stageD_evaluate_jump_target_add_29_U88 : XNOR2_X1 port map( A => 
                           n17178, B => 
                           pipeline_stageD_evaluate_jump_target_add_29_n207, ZN
                           => pipeline_stageD_evaluate_jump_target_N45);
   pipeline_stageD_evaluate_jump_target_add_29_U89 : AOI22_X1 port map( A1 => 
                           pipeline_nextPC_IFID_DEC_12_port, A2 => 
                           pipeline_stageD_offset_to_jump_temp_12_port, B1 => 
                           n17444, B2 => n17459, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n207);
   pipeline_stageD_evaluate_jump_target_add_29_U87 : XNOR2_X1 port map( A => 
                           pipeline_nextPC_IFID_DEC_13_port, B => 
                           pipeline_stageD_offset_to_jump_temp_13_port, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n203);
   pipeline_stageD_evaluate_jump_target_add_29_U81 : AOI22_X1 port map( A1 => 
                           pipeline_nextPC_IFID_DEC_14_port, A2 => 
                           pipeline_stageD_offset_to_jump_temp_14_port, B1 => 
                           n17445, B2 => n17460, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n201);
   pipeline_stageD_evaluate_jump_target_add_29_U79 : XNOR2_X1 port map( A => 
                           pipeline_nextPC_IFID_DEC_15_port, B => 
                           pipeline_stageD_offset_to_jump_temp_15_port, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n197);
   pipeline_stageD_evaluate_jump_target_add_29_U73 : AOI22_X1 port map( A1 => 
                           pipeline_nextPC_IFID_DEC_16_port, A2 => 
                           pipeline_stageD_offset_to_jump_temp_16_port, B1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n194, B2
                           => n17461, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n195);
   pipeline_stageD_evaluate_jump_target_add_29_U71 : XNOR2_X1 port map( A => 
                           pipeline_nextPC_IFID_DEC_17_port, B => 
                           pipeline_stageD_offset_to_jump_temp_17_port, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n191);
   pipeline_stageD_evaluate_jump_target_add_29_U65 : AOI22_X1 port map( A1 => 
                           pipeline_nextPC_IFID_DEC_18_port, A2 => 
                           pipeline_stageD_offset_to_jump_temp_18_port, B1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n188, B2
                           => n17462, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n189);
   pipeline_stageD_evaluate_jump_target_add_29_U63 : XNOR2_X1 port map( A => 
                           pipeline_nextPC_IFID_DEC_19_port, B => 
                           pipeline_stageD_offset_to_jump_temp_19_port, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n185);
   pipeline_stageD_evaluate_jump_target_add_29_U55 : AOI22_X1 port map( A1 => 
                           pipeline_nextPC_IFID_DEC_20_port, A2 => 
                           pipeline_stageD_offset_to_jump_temp_20_port, B1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n180, B2
                           => n17463, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n181);
   pipeline_stageD_evaluate_jump_target_add_29_U53 : XNOR2_X1 port map( A => 
                           pipeline_nextPC_IFID_DEC_21_port, B => 
                           pipeline_stageD_offset_to_jump_temp_21_port, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n177);
   pipeline_stageD_evaluate_jump_target_add_29_U47 : AOI22_X1 port map( A1 => 
                           pipeline_nextPC_IFID_DEC_22_port, A2 => 
                           pipeline_stageD_offset_to_jump_temp_22_port, B1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n174, B2
                           => n17464, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n175);
   pipeline_stageD_evaluate_jump_target_add_29_U45 : XNOR2_X1 port map( A => 
                           pipeline_nextPC_IFID_DEC_23_port, B => 
                           pipeline_stageD_offset_to_jump_temp_23_port, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n171);
   pipeline_stageD_evaluate_jump_target_add_29_U39 : AOI22_X1 port map( A1 => 
                           pipeline_nextPC_IFID_DEC_24_port, A2 => 
                           pipeline_stageD_offset_to_jump_temp_24_port, B1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n168, B2
                           => n17465, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n169);
   pipeline_stageD_evaluate_jump_target_add_29_U37 : XNOR2_X1 port map( A => 
                           pipeline_nextPC_IFID_DEC_25_port, B => 
                           pipeline_stageD_offset_to_jump_temp_30_port, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n165);
   pipeline_stageD_evaluate_jump_target_add_29_U31 : AOI22_X1 port map( A1 => 
                           pipeline_nextPC_IFID_DEC_26_port, A2 => 
                           pipeline_stageD_offset_to_jump_temp_30_port, B1 => 
                           n17200, B2 => n17466, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n163);
   pipeline_stageD_evaluate_jump_target_add_29_U29 : XNOR2_X1 port map( A => 
                           pipeline_nextPC_IFID_DEC_27_port, B => 
                           pipeline_stageD_offset_to_jump_temp_30_port, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n159);
   pipeline_stageD_evaluate_jump_target_add_29_U23 : AOI22_X1 port map( A1 => 
                           pipeline_nextPC_IFID_DEC_28_port, A2 => 
                           pipeline_stageD_offset_to_jump_temp_30_port, B1 => 
                           n17200, B2 => n17467, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n157);
   pipeline_stageD_evaluate_jump_target_add_29_U120 : XOR2_X1 port map( A => 
                           net175543, B => pipeline_nextPC_IFID_DEC_0_port, Z 
                           => pipeline_stageD_evaluate_jump_target_N33);
   pipeline_stageD_evaluate_jump_target_add_29_U119 : XOR2_X1 port map( A => 
                           pipeline_nextPC_IFID_DEC_1_port, B => 
                           pipeline_stageD_offset_to_jump_temp_1_port, Z => 
                           pipeline_stageD_evaluate_jump_target_add_29_n184);
   U10950 : NOR2_X1 port map( A1 => pipeline_inst_IFID_DEC_31_port, A2 => 
                           pipeline_inst_IFID_DEC_28_port, ZN => n14190);
   U10948 : NAND2_X1 port map( A1 => n14190, A2 => n17382, ZN => n14177);
   U10947 : NOR3_X1 port map( A1 => Rst, A2 => n17313, A3 => n14177, ZN => 
                           n13979);
   U11908 : INV_X1 port map( A => addr_to_dataRam_2_port, ZN => n17012);
   U11734 : NAND2_X1 port map( A1 => addr_to_dataRam_4_port, A2 => 
                           addr_to_dataRam_3_port, ZN => n17013);
   U11873 : INV_X1 port map( A => addr_to_dataRam_3_port, ZN => n17015);
   U11253 : OAI21_X2 port map( B1 => n17662, B2 => n17321, A => n16701, ZN => 
                           pipeline_stageE_input1_to_ALU_1_port);
   U8598 : NOR2_X2 port map( A1 => Rst, A2 => 
                           pipeline_WB_controls_in_MEMWB_0_port, ZN => n14134);
   U9351 : NOR2_X2 port map( A1 => n14860, A2 => n14866, ZN => n14223);
   U9340 : NOR2_X2 port map( A1 => n14865, A2 => n14861, ZN => n14214);
   U9337 : NOR2_X2 port map( A1 => n14863, A2 => n14861, ZN => n14212);
   U9334 : NOR2_X2 port map( A1 => n14860, A2 => n14861, ZN => n14210);
   U9343 : NOR2_X2 port map( A1 => n14864, A2 => n14861, ZN => n14216);
   U10234 : NOR3_X1 port map( A1 => n17409, A2 => n17313, A3 => n14177, ZN => 
                           n14947);
   U11803 : AND3_X2 port map( A1 => n17012, A2 => n17015, A3 => 
                           addr_to_dataRam_4_port, ZN => n16822);
   U10243 : NAND2_X1 port map( A1 => n17703, A2 => n15646, ZN => n14168);
   U10242 : INV_X1 port map( A => n14168, ZN => n14167);
   pipeline_stageF_PC_reg_PC_out_reg_30_inst : DFFR_X1 port map( D => n3989, CK
                           => Clk, RN => n17703, Q => n13782, QN => n7710);
   pipeline_IFID_stage_Instr_out_IFID_reg_1_inst : DFF_X2 port map( D => n3986,
                           CK => Clk, Q => 
                           pipeline_stageD_offset_to_jump_temp_1_port, QN => 
                           n17406);
   U12262 : OAI21_X1 port map( B1 => n14127, B2 => n17018, A => n17704, ZN => 
                           n14122);
   U12263 : OR2_X1 port map( A1 => n14125, A2 => n14126, ZN => n17018);
   U12264 : AOI222_X1 port map( A1 => n15598, A2 => n17579, B1 => n15598, B2 =>
                           pipeline_stageE_input1_to_ALU_3_port, C1 => n16688, 
                           C2 => pipeline_stageE_input1_to_ALU_3_port, ZN => 
                           n15566);
   U12265 : INV_X1 port map( A => pipeline_stageE_input1_to_ALU_30_port, ZN => 
                           n17083);
   U12266 : INV_X1 port map( A => pipeline_stageE_input1_to_ALU_19_port, ZN => 
                           n17097);
   U12267 : INV_X1 port map( A => pipeline_stageE_input1_to_ALU_5_port, ZN => 
                           n17087);
   U12268 : AND2_X1 port map( A1 => n17019, A2 => n17020, ZN => n12766);
   U12269 : BUF_X2 port map( A => n12766, Z => n17155);
   U12270 : NOR2_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_0_port, A2
                           => n13846, ZN => n17021);
   U12271 : AOI22_X1 port map( A1 => n17666, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_3_port, B1 => 
                           pipeline_data_to_RF_from_WB_3_port, B2 => n15123, ZN
                           => n17022);
   U12272 : OAI21_X1 port map( B1 => n17642, B2 => n17021, A => n17022, ZN => 
                           n17023);
   U12273 : OAI21_X2 port map( B1 => pipeline_immediate_to_exe_3_port, B2 => 
                           n17327, A => n17023, ZN => n17739);
   U12274 : NAND4_X1 port map( A1 => n15045, A2 => n14970, A3 => n14948, A4 => 
                           n15046, ZN => n17024);
   U12275 : NOR4_X1 port map( A1 => n15041, A2 => n15042, A3 => n15043, A4 => 
                           n17024, ZN => n17025);
   U12276 : NAND2_X1 port map( A1 => n17025, A2 => n15037, ZN => n17026);
   U12277 : NOR4_X1 port map( A1 => n15035, A2 => n15033, A3 => n15034, A4 => 
                           n17026, ZN => n17027);
   U12278 : AND4_X1 port map( A1 => n15039, A2 => n15040, A3 => n17027, A4 => 
                           n15032, ZN => n17028);
   U12279 : NAND3_X1 port map( A1 => n15030, A2 => n15029, A3 => n17028, ZN => 
                           n17029);
   U12280 : NOR4_X1 port map( A1 => n15026, A2 => n15025, A3 => n15027, A4 => 
                           n17029, ZN => n17030);
   U12281 : NAND2_X1 port map( A1 => n15017, A2 => n17030, ZN => n17538);
   U12282 : AOI21_X1 port map( B1 => n15138, B2 => n15137, A => n17608, ZN => 
                           n17031);
   U12283 : AOI21_X1 port map( B1 => n15142, B2 => n17542, A => n17031, ZN => 
                           n17032);
   U12284 : AOI21_X1 port map( B1 => n17104, B2 => n15137, A => n17032, ZN => 
                           n15005);
   U12285 : OR2_X1 port map( A1 => n17327, A2 => 
                           pipeline_immediate_to_exe_1_port, ZN => n17033);
   U12286 : OAI21_X1 port map( B1 => n17642, B2 => n17577, A => n16699, ZN => 
                           n17034);
   U12287 : NAND2_X1 port map( A1 => n17034, A2 => n17033, ZN => n17741);
   U12288 : NOR4_X1 port map( A1 => n15022, A2 => n15021, A3 => n15023, A4 => 
                           n15024, ZN => n17035);
   U12289 : NAND2_X1 port map( A1 => n15020, A2 => n17035, ZN => n17537);
   U12290 : INV_X1 port map( A => n17411, ZN => n17036);
   U12291 : NOR3_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_2_port, A2
                           => pipeline_EXE_controls_in_EXEcute_4_port, A3 => 
                           n17036, ZN => n17528);
   U12292 : AOI22_X1 port map( A1 => n17742, A2 => 
                           pipeline_stageE_EXE_ALU_add_alu_sCout_0_port, B1 => 
                           pipeline_stageE_input2_to_ALU_0_port, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N202, ZN => n15048
                           );
   U12293 : AOI22_X1 port map( A1 => n17664, A2 => n13832, B1 => n17663, B2 => 
                           pipeline_Alu_Out_Addr_to_mem_5_port, ZN => n17037);
   U12294 : OAI21_X1 port map( B1 => n17105, B2 => n17308, A => n17037, ZN => 
                           pipeline_stageE_input1_to_ALU_5_port);
   U12295 : NOR2_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_0_port, A2
                           => n13811, ZN => n17038);
   U12296 : OAI21_X1 port map( B1 => n17642, B2 => n17038, A => n16704, ZN => 
                           n17039);
   U12297 : OAI21_X1 port map( B1 => pipeline_immediate_to_exe_2_port, B2 => 
                           n17327, A => n17039, ZN => n17740);
   U12298 : OAI21_X1 port map( B1 => n17166, B2 => 
                           pipeline_stageD_offset_to_jump_temp_23_port, A => 
                           pipeline_nextPC_IFID_DEC_23_port, ZN => n17196);
   U12299 : AOI222_X1 port map( A1 => pipeline_Alu_Out_Addr_to_mem_30_port, A2 
                           => n17331, B1 => n13782, B2 => n17674, C1 => n17108,
                           C2 => pipeline_stageF_PC_plus4_N37, ZN => n17638);
   U12300 : AND3_X1 port map( A1 => n15383, A2 => n15368, A3 => n15367, ZN => 
                           n17040);
   U12301 : NOR2_X1 port map( A1 => n17040, A2 => n15352, ZN => n17041);
   U12302 : XNOR2_X1 port map( A => n17041, B => n17096, ZN => n17042);
   U12303 : XNOR2_X1 port map( A => n17042, B => n15348, ZN => n15021);
   U12304 : INV_X1 port map( A => n17121, ZN => n17043);
   U12305 : AOI222_X1 port map( A1 => n17043, A2 => 
                           pipeline_data_to_RF_from_WB_2_port, B1 => n17663, B2
                           => pipeline_Alu_Out_Addr_to_mem_2_port, C1 => n16620
                           , C2 => n13809, ZN => n17044);
   U12306 : INV_X1 port map( A => n17044, ZN => n12649);
   U12307 : AOI22_X1 port map( A1 => n17428, A2 => n17457, B1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n128, B2
                           => n17295, ZN => n17177);
   U12308 : NOR4_X1 port map( A1 => n16554, A2 => n16796, A3 => n16795, A4 => 
                           n17387, ZN => n16619);
   U12309 : NAND2_X1 port map( A1 => pipeline_stageE_input1_to_ALU_23_port, A2 
                           => n15263, ZN => n17045);
   U12310 : AOI21_X1 port map( B1 => n15265, B2 => n17045, A => n17603, ZN => 
                           n17046);
   U12311 : NAND2_X1 port map( A1 => n17045, A2 => n15268, ZN => n17047);
   U12312 : OAI21_X1 port map( B1 => n15282, B2 => n17047, A => n17046, ZN => 
                           n15248);
   U12313 : AOI22_X1 port map( A1 => n17739, A2 => n17381, B1 => 
                           pipeline_stageE_EXE_ALU_add_alu_sCout_0_port, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_3_port, ZN 
                           => n15598);
   U12314 : NAND4_X1 port map( A1 => n17279, A2 => n17278, A3 => 
                           pipeline_nextPC_IFID_DEC_29_port, A4 => n17183, ZN 
                           => n17186);
   U12315 : AOI222_X1 port map( A1 => n15368, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_A_16_port, B1 
                           => n15368, B2 => n15369, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_A_16_port, C2 
                           => n15369, ZN => n17048);
   U12316 : NAND2_X1 port map( A1 => n15367, A2 => n15366, ZN => n17049);
   U12317 : XOR2_X1 port map( A => n17048, B => n17049, Z => n15025);
   U12318 : INV_X1 port map( A => n14094, ZN => n17050);
   U12319 : AOI22_X1 port map( A1 => n14094, A2 => 
                           pipeline_stageD_offset_jump_sign_ext_24_port, B1 => 
                           pipeline_stageD_offset_jump_sign_ext_19_port, B2 => 
                           n17050, ZN => n17051);
   U12320 : AOI22_X1 port map( A1 => n14094, A2 => 
                           pipeline_stageD_offset_jump_sign_ext_31_port, B1 => 
                           pipeline_stageD_offset_jump_sign_ext_20_port, B2 => 
                           n17050, ZN => n17052);
   U12321 : NOR3_X1 port map( A1 => n14091, A2 => n14087, A3 => n14098, ZN => 
                           n17053);
   U12322 : OAI22_X1 port map( A1 => n14116, A2 => 
                           pipeline_stageD_offset_jump_sign_ext_16_port, B1 => 
                           pipeline_stageD_offset_jump_sign_ext_17_port, B2 => 
                           n14117, ZN => n17054);
   U12323 : AOI221_X1 port map( B1 => n14116, B2 => 
                           pipeline_stageD_offset_jump_sign_ext_16_port, C1 => 
                           n14117, C2 => 
                           pipeline_stageD_offset_jump_sign_ext_17_port, A => 
                           n17054, ZN => n17055);
   U12324 : OAI211_X1 port map( C1 => n14113, C2 => 
                           pipeline_stageD_offset_jump_sign_ext_18_port, A => 
                           n17055, B => n14091, ZN => n17056);
   U12325 : AOI21_X1 port map( B1 => n14113, B2 => 
                           pipeline_stageD_offset_jump_sign_ext_18_port, A => 
                           n17056, ZN => n17057);
   U12326 : XNOR2_X1 port map( A => n14101, B => n17052, ZN => n17058);
   U12327 : OAI21_X1 port map( B1 => n17057, B2 => n17053, A => n17058, ZN => 
                           n17059);
   U12328 : XOR2_X1 port map( A => n14100, B => n17051, Z => n17060);
   U12329 : NOR3_X1 port map( A1 => n17060, A2 => n14096, A3 => n17059, ZN => 
                           n14092);
   U12330 : NAND4_X1 port map( A1 => pipeline_inst_IFID_DEC_29_port, A2 => 
                           n14049, A3 => n13993, A4 => 
                           pipeline_inst_IFID_DEC_27_port, ZN => n17061);
   U12331 : OAI211_X1 port map( C1 => n14059, C2 => n14058, A => n14020, B => 
                           n17061, ZN => n17062);
   U12332 : NOR2_X1 port map( A1 => n17350, A2 => n14064, ZN => n17063);
   U12333 : AOI21_X1 port map( B1 => n14065, B2 => n17076, A => n17063, ZN => 
                           n17064);
   U12334 : AOI221_X1 port map( B1 => n14066, B2 => n17064, C1 => n17076, C2 =>
                           n17064, A => n14012, ZN => n17065);
   U12335 : AOI211_X1 port map( C1 => n14032, C2 => n14033, A => n17062, B => 
                           n17065, ZN => n14041);
   U12336 : OAI221_X1 port map( B1 => n15000, B2 => 
                           pipeline_EXE_controls_in_EXEcute_2_port, C1 => 
                           n15000, C2 => n15001, A => n17529, ZN => n17066);
   U12337 : AOI21_X1 port map( B1 => n14964, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N105, A => n17623,
                           ZN => n17067);
   U12338 : NAND2_X1 port map( A1 => n17066, A2 => n17067, ZN => 
                           pipeline_EXMEM_stage_N7);
   U12339 : INV_X1 port map( A => n17106, ZN => n17068);
   U12340 : NAND2_X1 port map( A1 => n17330, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_29_port, ZN => n17069);
   U12341 : NAND3_X1 port map( A1 => n17069, A2 => n17622, A3 => n17621, ZN => 
                           n17070);
   U12342 : AOI21_X1 port map( B1 => pipeline_data_to_RF_from_WB_29_port, B2 =>
                           n17332, A => n17070, ZN => n17071);
   U12343 : NAND2_X1 port map( A1 => n15607, A2 => 
                           pipeline_stageD_target_Jump_temp_29_port, ZN => 
                           n17072);
   U12344 : OAI211_X1 port map( C1 => n14887, C2 => n17068, A => n17071, B => 
                           n17072, ZN => n3988);
   U12345 : AND2_X2 port map( A1 => n17233, A2 => n17232, ZN => n17162);
   U12346 : AND2_X2 port map( A1 => n17263, A2 => n17262, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n133);
   U12347 : INV_X1 port map( A => n17740, ZN => n17073);
   U12348 : INV_X4 port map( A => n17740, ZN => n17074);
   U12349 : NOR2_X2 port map( A1 => n16691, A2 => n12649, ZN => n15055);
   U12350 : NAND2_X4 port map( A1 => n14025, A2 => n14167, ZN => n17075);
   U12351 : INV_X2 port map( A => n4376, ZN => n17737);
   U12352 : NOR2_X4 port map( A1 => n15648, A2 => n15646, ZN => n15600);
   U12353 : BUF_X4 port map( A => pipeline_stageE_EXE_ALU_alu_shift_C86_n27, Z 
                           => n17111);
   U12354 : OAI21_X2 port map( B1 => n17662, B2 => n17306, A => n16689, ZN => 
                           pipeline_stageE_input1_to_ALU_3_port);
   U12355 : INV_X2 port map( A => pipeline_stageE_input2_to_ALU_0_port, ZN => 
                           n17742);
   U12356 : NOR2_X2 port map( A1 => n17387, A2 => n14982, ZN => n16607);
   U12357 : INV_X2 port map( A => n17741, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_1_port);
   U12358 : INV_X4 port map( A => n17302, ZN => n17112);
   U12359 : INV_X4 port map( A => n17303, ZN => n17099);
   U12360 : CLKBUF_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_3_port, Z 
                           => n17300);
   U12361 : CLKBUF_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_3_port, Z 
                           => n17301);
   U12362 : CLKBUF_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_3_port, Z 
                           => n17299);
   U12363 : CLKBUF_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_1_port, Z 
                           => n17298);
   U12364 : INV_X2 port map( A => n17739, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_3_port);
   U12365 : INV_X2 port map( A => Rst, ZN => n17703);
   U12366 : AOI21_X1 port map( B1 => n17164, B2 => 
                           pipeline_nextPC_IFID_DEC_25_port, A => n17202, ZN =>
                           pipeline_stageD_evaluate_jump_target_add_29_n160);
   U12367 : AOI222_X2 port map( A1 => pipeline_nextPC_IFID_DEC_1_port, A2 => 
                           pipeline_stageD_offset_to_jump_temp_1_port, B1 => 
                           n17167, B2 => pipeline_nextPC_IFID_DEC_1_port, C1 =>
                           pipeline_stageD_evaluate_jump_target_add_29_n214, C2
                           => pipeline_stageD_offset_to_jump_temp_1_port, ZN =>
                           n17161);
   U12368 : INV_X1 port map( A => pipeline_stageE_EXE_ALU_alu_shift_N136, ZN =>
                           n17104);
   U12369 : INV_X1 port map( A => pipeline_stageE_input1_to_ALU_3_port, ZN => 
                           n17077);
   U12370 : INV_X1 port map( A => pipeline_stageE_input1_to_ALU_27_port, ZN => 
                           n17078);
   U12371 : INV_X1 port map( A => pipeline_stageE_input1_to_ALU_17_port, ZN => 
                           n17079);
   U12372 : INV_X1 port map( A => pipeline_stageE_input1_to_ALU_12_port, ZN => 
                           n17080);
   U12373 : INV_X1 port map( A => n17074, ZN => n17081);
   U12374 : INV_X1 port map( A => pipeline_stageE_input1_to_ALU_11_port, ZN => 
                           n17082);
   U12375 : INV_X1 port map( A => pipeline_stageE_input1_to_ALU_21_port, ZN => 
                           n17084);
   U12376 : INV_X1 port map( A => pipeline_stageE_input1_to_ALU_10_port, ZN => 
                           n17085);
   U12377 : OAI21_X1 port map( B1 => n17121, B2 => n17320, A => n16684, ZN => 
                           pipeline_stageE_input1_to_ALU_4_port);
   U12378 : INV_X1 port map( A => pipeline_stageE_input1_to_ALU_26_port, ZN => 
                           n17086);
   U12379 : INV_X1 port map( A => pipeline_stageE_input1_to_ALU_6_port, ZN => 
                           n17088);
   U12380 : INV_X1 port map( A => pipeline_stageE_input1_to_ALU_7_port, ZN => 
                           n17089);
   U12381 : INV_X1 port map( A => pipeline_stageE_input1_to_ALU_9_port, ZN => 
                           n17090);
   U12382 : INV_X1 port map( A => n12649, ZN => n17091);
   U12383 : INV_X1 port map( A => pipeline_stageE_input1_to_ALU_23_port, ZN => 
                           n17092);
   U12384 : INV_X1 port map( A => pipeline_stageE_input1_to_ALU_28_port, ZN => 
                           n17093);
   U12385 : INV_X1 port map( A => pipeline_stageE_input1_to_ALU_29_port, ZN => 
                           n17094);
   U12386 : INV_X1 port map( A => pipeline_stageE_input1_to_ALU_8_port, ZN => 
                           n17095);
   U12387 : INV_X1 port map( A => pipeline_stageE_input1_to_ALU_18_port, ZN => 
                           n17096);
   U12388 : NAND2_X2 port map( A1 => n17703, A2 => n17422, ZN => n17418);
   U12389 : BUF_X1 port map( A => n16591, Z => n17658);
   U12390 : BUF_X1 port map( A => n16595, Z => n17654);
   U12391 : BUF_X1 port map( A => n13151, Z => n17713);
   U12392 : INV_X2 port map( A => n16777, ZN => n17120);
   U12393 : AND2_X1 port map( A1 => n17572, A2 => n17662, ZN => n16620);
   U12394 : BUF_X1 port map( A => n16592, Z => n17657);
   U12395 : BUF_X1 port map( A => n16593, Z => n17656);
   U12396 : BUF_X1 port map( A => n16594, Z => n17655);
   U12397 : BUF_X1 port map( A => n16596, Z => n17651);
   U12398 : BUF_X1 port map( A => n16597, Z => n17650);
   U12399 : BUF_X1 port map( A => n16590, Z => n17661);
   U12400 : NAND2_X2 port map( A1 => n17670, A2 => n13942, ZN => n17422);
   U12401 : BUF_X1 port map( A => n16617, Z => n17105);
   U12402 : NOR2_X1 port map( A1 => n17012, A2 => n17013, ZN => n17660);
   U12403 : NOR2_X2 port map( A1 => addr_to_dataRam_2_port, A2 => n17013, ZN =>
                           n17530);
   U12404 : BUF_X2 port map( A => n13055, Z => n17098);
   U12405 : BUF_X1 port map( A => n17672, Z => n17107);
   U12406 : NOR2_X1 port map( A1 => pipeline_stall, A2 => n15648, ZN => n17672)
                           ;
   U12407 : INV_X1 port map( A => n17420, ZN => n17109);
   U12408 : AOI221_X1 port map( B1 => pipeline_stageE_EXE_ALU_alu_shift_C50_n51
                           , B2 => pipeline_stageE_input1_to_ALU_14_port, C1 =>
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n167, C2 => 
                           n17160, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n132, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n43);
   U12409 : AOI221_X1 port map( B1 => pipeline_stageE_EXE_ALU_alu_shift_C48_n2,
                           B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_A_16_port, C1 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_n53, C2 => 
                           pipeline_stageE_input1_to_ALU_17_port, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n151, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n115);
   U12410 : AOI221_X1 port map( B1 => pipeline_stageE_EXE_ALU_alu_shift_C50_n51
                           , B2 => n17160, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n167, C2 => 
                           pipeline_stageE_input1_to_ALU_12_port, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n144, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n63);
   U12411 : AOI221_X1 port map( B1 => pipeline_stageE_EXE_ALU_alu_shift_C48_n2,
                           B2 => pipeline_stageE_input1_to_ALU_14_port, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n53, C2 => 
                           pipeline_stageE_input1_to_ALU_15_port, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n161, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n134);
   U12412 : AOI221_X1 port map( B1 => n17156, B2 => 
                           pipeline_stageE_input1_to_ALU_6_port, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n53, C2 => 
                           pipeline_stageE_input1_to_ALU_7_port, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n170, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n36);
   U12413 : AOI221_X1 port map( B1 => n17156, B2 => 
                           pipeline_stageE_input1_to_ALU_7_port, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n53, C2 => 
                           pipeline_stageE_input1_to_ALU_8_port, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n100, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n32);
   U12414 : AOI221_X1 port map( B1 => pipeline_stageE_EXE_ALU_alu_shift_C48_n2,
                           B2 => pipeline_stageE_input1_to_ALU_8_port, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n53, C2 => 
                           pipeline_stageE_input1_to_ALU_9_port, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n67, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n26);
   U12415 : AOI221_X1 port map( B1 => n17156, B2 => 
                           pipeline_stageE_input1_to_ALU_9_port, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n53, C2 => 
                           pipeline_stageE_input1_to_ALU_10_port, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n54, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n20);
   U12416 : INV_X2 port map( A => pipeline_stall, ZN => n15646);
   U12417 : NAND2_X1 port map( A1 => n16693, A2 => 
                           pipeline_stageE_input1_to_ALU_1_port, ZN => n15049);
   U12418 : NAND2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_1_port, A2 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, 
                           ZN => pipeline_stageE_EXE_ALU_alu_shift_C50_n44);
   U12419 : OAI21_X1 port map( B1 => n17121, B2 => n17362, A => n16792, ZN => 
                           pipeline_stageE_input1_to_ALU_30_port);
   U12420 : INV_X1 port map( A => pipeline_stageE_input1_to_ALU_14_port, ZN => 
                           n17100);
   U12421 : INV_X1 port map( A => pipeline_stageE_input1_to_ALU_15_port, ZN => 
                           n17101);
   U12422 : INV_X1 port map( A => pipeline_stageE_input1_to_ALU_4_port, ZN => 
                           n17102);
   U12423 : INV_X1 port map( A => pipeline_stageE_input1_to_ALU_1_port, ZN => 
                           n17103);
   U12424 : NAND2_X1 port map( A1 => n17653, A2 => n17098, ZN => n16595);
   U12425 : BUF_X1 port map( A => n16617, Z => n17121);
   U12426 : BUF_X1 port map( A => n17652, Z => n17653);
   U12427 : BUF_X1 port map( A => n17668, Z => n17123);
   U12428 : NOR2_X1 port map( A1 => n17012, A2 => n17013, ZN => n16823);
   U12429 : BUF_X1 port map( A => n16817, Z => n17124);
   U12430 : NOR2_X2 port map( A1 => addr_to_dataRam_2_port, A2 => n17013, ZN =>
                           n16824);
   U12431 : NOR2_X1 port map( A1 => addr_to_dataRam_4_port, A2 => n17016, ZN =>
                           n16819);
   U12432 : BUF_X1 port map( A => n16818, Z => n17125);
   U12433 : NOR2_X1 port map( A1 => n17012, A2 => n17013, ZN => n17659);
   U12434 : INV_X1 port map( A => n16561, ZN => n17643);
   U12435 : BUF_X1 port map( A => n14964, Z => n17126);
   U12436 : NOR2_X2 port map( A1 => addr_to_dataRam_3_port, A2 => n17014, ZN =>
                           n17531);
   U12437 : NOR2_X1 port map( A1 => n17155, A2 => read_notWrite, ZN => n13055);
   U12438 : NOR2_X2 port map( A1 => addr_to_dataRam_3_port, A2 => n17014, ZN =>
                           n16821);
   U12439 : NOR2_X2 port map( A1 => pipeline_EXE_controls_in_EXEcute_3_port, A2
                           => n15582, ZN => n17419);
   U12440 : BUF_X1 port map( A => n15903, Z => n17142);
   U12441 : BUF_X1 port map( A => n15931, Z => n17145);
   U12442 : BUF_X1 port map( A => n15918, Z => n17141);
   U12443 : BUF_X1 port map( A => n15905, Z => n17144);
   U12444 : BUF_X1 port map( A => n15914, Z => n17136);
   U12445 : BUF_X1 port map( A => n15912, Z => n17140);
   U12446 : BUF_X1 port map( A => n15930, Z => n17143);
   U12447 : BUF_X1 port map( A => n15917, Z => n17139);
   U12448 : BUF_X1 port map( A => n15926, Z => n17148);
   U12449 : BUF_X1 port map( A => n15927, Z => n17131);
   U12450 : BUF_X1 port map( A => n15924, Z => n17128);
   U12451 : BUF_X1 port map( A => n15928, Z => n17146);
   U12452 : BUF_X1 port map( A => n15925, Z => n17134);
   U12453 : BUF_X1 port map( A => n15929, Z => n17147);
   U12454 : BUF_X1 port map( A => n15940, Z => n17137);
   U12455 : BUF_X1 port map( A => n15935, Z => n17135);
   U12456 : BUF_X1 port map( A => n15936, Z => n17132);
   U12457 : BUF_X1 port map( A => n15937, Z => n17127);
   U12458 : BUF_X1 port map( A => n15906, Z => n17133);
   U12459 : BUF_X1 port map( A => n15941, Z => n17138);
   U12460 : BUF_X1 port map( A => n15938, Z => n17130);
   U12461 : BUF_X1 port map( A => n15939, Z => n17129);
   U12462 : NOR2_X2 port map( A1 => n14860, A2 => n14866, ZN => n17417);
   U12463 : NOR2_X2 port map( A1 => n14864, A2 => n14861, ZN => n17413);
   U12464 : NOR2_X2 port map( A1 => n14865, A2 => n14861, ZN => n17414);
   U12465 : NOR2_X2 port map( A1 => n14863, A2 => n14861, ZN => n17415);
   U12466 : NOR2_X2 port map( A1 => n14860, A2 => n14861, ZN => n17416);
   U12467 : AOI221_X1 port map( B1 => n17304, B2 => 
                           pipeline_stageD_offset_jump_sign_ext_22_port, C1 => 
                           pipeline_stageD_offset_jump_sign_ext_31_port, C2 => 
                           n17386, A => n16568, ZN => n16565);
   U12468 : NOR2_X2 port map( A1 => Rst, A2 => 
                           pipeline_WB_controls_in_MEMWB_0_port, ZN => n17370);
   U12469 : INV_X1 port map( A => Rst, ZN => n17701);
   U12470 : INV_X1 port map( A => Rst, ZN => n17702);
   U12471 : INV_X2 port map( A => Rst, ZN => n17704);
   U12472 : NOR3_X1 port map( A1 => n17606, A2 => n17605, A3 => n17604, ZN => 
                           n15218);
   U12473 : AOI21_X1 port map( B1 => n16646, B2 => n17591, A => n17592, ZN => 
                           n15368);
   U12474 : AND3_X1 port map( A1 => n17588, A2 => n17589, A3 => n17590, ZN => 
                           n15445);
   U12475 : BUF_X1 port map( A => n15600, Z => n17671);
   U12476 : BUF_X1 port map( A => n15601, Z => n17673);
   U12477 : BUF_X2 port map( A => n15608, Z => n17106);
   U12478 : BUF_X2 port map( A => n15610, Z => n17108);
   U12479 : AOI221_X1 port map( B1 => pipeline_stageE_EXE_ALU_alu_shift_C48_n2,
                           B2 => pipeline_stageE_input1_to_ALU_15_port, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n53, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_A_16_port, A 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_n132, ZN =>
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n99);
   U12480 : BUF_X1 port map( A => n15611, Z => n17674);
   U12481 : AOI221_X1 port map( B1 => pipeline_stageE_EXE_ALU_alu_shift_C48_n2,
                           B2 => pipeline_stageE_input1_to_ALU_11_port, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n53, C2 => 
                           pipeline_stageE_input1_to_ALU_12_port, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n94, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n4);
   U12482 : AOI221_X1 port map( B1 => pipeline_stageE_EXE_ALU_alu_shift_C48_n2,
                           B2 => pipeline_stageE_input1_to_ALU_13_port, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n53, C2 => 
                           pipeline_stageE_input1_to_ALU_14_port, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n145, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n45);
   U12483 : AOI221_X1 port map( B1 => pipeline_stageE_EXE_ALU_alu_shift_C48_n2,
                           B2 => pipeline_stageE_input1_to_ALU_12_port, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n53, C2 => 
                           n17160, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n154, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n64);
   U12484 : AOI221_X1 port map( B1 => pipeline_stageE_EXE_ALU_alu_shift_C48_n2,
                           B2 => pipeline_stageE_input1_to_ALU_10_port, C1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n53, C2 => 
                           pipeline_stageE_input1_to_ALU_11_port, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n157, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n14);
   U12485 : BUF_X2 port map( A => pipeline_stageE_EXE_ALU_alu_shift_C86_n26, Z 
                           => n17110);
   U12486 : NAND2_X2 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_1_port, A2 
                           => n17742, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n21);
   U12487 : NAND2_X2 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, A2 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_SH_1_port, 
                           ZN => pipeline_stageE_EXE_ALU_alu_shift_C86_n23);
   U12488 : BUF_X2 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, Z 
                           => n17113);
   U12489 : INV_X2 port map( A => n17081, ZN => n17114);
   U12490 : INV_X1 port map( A => pipeline_stageE_input1_to_ALU_25_port, ZN => 
                           n17115);
   U12491 : INV_X1 port map( A => pipeline_stageE_input1_to_ALU_22_port, ZN => 
                           n17116);
   U12492 : INV_X1 port map( A => pipeline_stageE_input1_to_ALU_24_port, ZN => 
                           n17117);
   U12493 : INV_X1 port map( A => pipeline_stageE_input1_to_ALU_20_port, ZN => 
                           n17118);
   U12494 : INV_X1 port map( A => pipeline_stageE_EXE_ALU_alu_shift_N202, ZN =>
                           n17119);
   U12495 : BUF_X1 port map( A => n16620, Z => n17664);
   U12496 : BUF_X1 port map( A => n13103, Z => n17729);
   U12497 : NAND2_X1 port map( A1 => n17530, A2 => n17098, ZN => n16591);
   U12498 : BUF_X1 port map( A => n16617, Z => n17662);
   U12499 : BUF_X1 port map( A => n17669, Z => n17670);
   U12500 : BUF_X2 port map( A => n16619, Z => n17663);
   U12501 : BUF_X2 port map( A => n16819, Z => n17122);
   U12502 : NOR3_X1 port map( A1 => addr_to_dataRam_4_port, A2 => 
                           addr_to_dataRam_2_port, A3 => n17015, ZN => n17652);
   U12503 : NAND2_X2 port map( A1 => 
                           pipeline_stageE_EXE_ALU_add_alu_sCout_0_port, A2 => 
                           n15573, ZN => n14968);
   U12504 : BUF_X2 port map( A => n14213, Z => n17700);
   U12505 : BUF_X1 port map( A => n14246, Z => n17687);
   U12506 : BUF_X2 port map( A => n14225, Z => n17698);
   U12507 : BUF_X1 port map( A => n14238, Z => n17691);
   U12508 : BUF_X1 port map( A => n14250, Z => n17683);
   U12509 : BUF_X1 port map( A => n14240, Z => n17689);
   U12510 : BUF_X2 port map( A => n14247, Z => n17684);
   U12511 : BUF_X2 port map( A => n14239, Z => n17688);
   U12512 : BUF_X1 port map( A => n14248, Z => n17685);
   U12513 : BUF_X1 port map( A => n14222, Z => n17699);
   U12514 : BUF_X2 port map( A => n14244, Z => n17686);
   U12515 : BUF_X1 port map( A => n14236, Z => n17693);
   U12516 : BUF_X1 port map( A => n14234, Z => n17695);
   U12517 : BUF_X2 port map( A => n14227, Z => n17696);
   U12518 : BUF_X2 port map( A => n14237, Z => n17690);
   U12519 : BUF_X1 port map( A => n14228, Z => n17697);
   U12520 : BUF_X2 port map( A => n14233, Z => n17694);
   U12521 : BUF_X2 port map( A => n14235, Z => n17692);
   U12522 : NOR2_X2 port map( A1 => n16529, A2 => n16531, ZN => n17392);
   U12523 : NOR2_X2 port map( A1 => n16530, A2 => n16534, ZN => n17390);
   U12524 : NOR2_X2 port map( A1 => n16532, A2 => n16534, ZN => n17389);
   U12525 : NOR2_X2 port map( A1 => n16527, A2 => n16534, ZN => n17388);
   U12526 : NOR2_X2 port map( A1 => n16527, A2 => n16528, ZN => n17391);
   U12527 : BUF_X2 port map( A => n14966, Z => n17149);
   U12528 : BUF_X2 port map( A => n14965, Z => n17150);
   U12529 : BUF_X2 port map( A => n14215, Z => n17151);
   U12530 : BUF_X2 port map( A => n14224, Z => n17152);
   U12531 : BUF_X2 port map( A => n14245, Z => n17153);
   U12532 : BUF_X2 port map( A => n14249, Z => n17154);
   U12533 : CLKBUF_X1 port map( A => pipeline_Forward_sw1_mux, Z => n17744);
   U12534 : INV_X1 port map( A => pipeline_Forward_sw1_mux, ZN => n17743);
   U12535 : NOR2_X2 port map( A1 => n16530, A2 => n16534, ZN => n15913);
   U12536 : NOR2_X2 port map( A1 => n16532, A2 => n16534, ZN => n15915);
   U12537 : NOR2_X2 port map( A1 => n16527, A2 => n16528, ZN => n15901);
   U12538 : NOR2_X2 port map( A1 => pipeline_EXE_controls_in_EXEcute_3_port, A2
                           => n15582, ZN => n14961);
   U12539 : OAI21_X2 port map( B1 => n17105, B2 => n17425, A => n16793, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N136);
   U12540 : INV_X1 port map( A => pipeline_stageE_EXE_ALU_alu_shift_C48_n46, ZN
                           => n17156);
   U12541 : NOR2_X2 port map( A1 => n17742, A2 => n17303, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n53);
   U12542 : NOR2_X2 port map( A1 => n17411, A2 => n15588, ZN => n14954);
   U12543 : INV_X1 port map( A => n17118, ZN => n17157);
   U12544 : NOR2_X2 port map( A1 => n17074, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_3_port, ZN 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_n1);
   U12545 : OAI21_X2 port map( B1 => n17662, B2 => n17318, A => n16678, ZN => 
                           pipeline_stageE_input1_to_ALU_6_port);
   U12546 : OAI21_X2 port map( B1 => n17121, B2 => n17423, A => n16637, ZN => 
                           pipeline_stageE_input1_to_ALU_19_port);
   U12547 : OAI21_X2 port map( B1 => n17105, B2 => n17363, A => n16734, ZN => 
                           pipeline_stageE_input1_to_ALU_18_port);
   U12548 : OAI21_X2 port map( B1 => n17105, B2 => n17365, A => n16770, ZN => 
                           pipeline_stageE_input1_to_ALU_29_port);
   U12549 : INV_X2 port map( A => n14981, ZN => n14952);
   U12550 : INV_X1 port map( A => n17117, ZN => n17158);
   U12551 : OAI21_X2 port map( B1 => n17105, B2 => n17309, A => n16653, ZN => 
                           pipeline_stageE_input1_to_ALU_14_port);
   U12552 : OAI21_X2 port map( B1 => n17105, B2 => n17325, A => n16762, ZN => 
                           pipeline_stageE_input1_to_ALU_27_port);
   U12553 : OAI21_X2 port map( B1 => n17121, B2 => n17424, A => n16758, ZN => 
                           pipeline_stageE_input1_to_ALU_26_port);
   U12554 : OAI21_X2 port map( B1 => n17121, B2 => n17364, A => n16733, ZN => 
                           pipeline_stageE_input1_to_ALU_15_port);
   U12555 : OAI21_X2 port map( B1 => n17121, B2 => n17307, A => n16721, ZN => 
                           pipeline_stageE_input1_to_ALU_10_port);
   U12556 : OAI21_X2 port map( B1 => n17105, B2 => n17305, A => n16671, ZN => 
                           pipeline_stageE_input1_to_ALU_9_port);
   U12557 : INV_X1 port map( A => n17115, ZN => n17159);
   U12558 : OAI21_X2 port map( B1 => n17105, B2 => n17312, A => n16766, ZN => 
                           pipeline_stageE_input1_to_ALU_28_port);
   U12559 : OAI21_X2 port map( B1 => n17121, B2 => n17343, A => n16713, ZN => 
                           pipeline_stageE_input1_to_ALU_7_port);
   U12560 : OAI21_X2 port map( B1 => n17121, B2 => n17394, A => n16720, ZN => 
                           pipeline_stageE_input1_to_ALU_8_port);
   U12561 : OAI21_X2 port map( B1 => n17121, B2 => n17395, A => n16660, ZN => 
                           pipeline_stageE_input1_to_ALU_12_port);
   U12562 : OAI21_X2 port map( B1 => n17105, B2 => n17323, A => n16645, ZN => 
                           pipeline_stageE_input1_to_ALU_17_port);
   U12563 : OAI21_X2 port map( B1 => n17105, B2 => n17319, A => n16725, ZN => 
                           pipeline_stageE_input1_to_ALU_11_port);
   U12564 : OAI21_X2 port map( B1 => n17121, B2 => n17311, A => n16749, ZN => 
                           pipeline_stageE_input1_to_ALU_22_port);
   U12565 : OAI21_X2 port map( B1 => n17121, B2 => n17310, A => n16742, ZN => 
                           pipeline_stageE_input1_to_ALU_21_port);
   U12566 : OAI21_X2 port map( B1 => n17105, B2 => n17366, A => n16753, ZN => 
                           pipeline_stageE_input1_to_ALU_23_port);
   U12567 : INV_X1 port map( A => n15425, ZN => n17160);
   U12568 : INV_X4 port map( A => n17742, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port);
   U12569 : NOR4_X2 port map( A1 => pipeline_stageD_offset_to_jump_temp_10_port
                           , A2 => pipeline_stageD_offset_to_jump_temp_9_port, 
                           A3 => pipeline_stageD_offset_to_jump_temp_7_port, A4
                           => n14174, ZN => n14005);
   U12570 : NOR2_X2 port map( A1 => n16529, A2 => n16531, ZN => n15907);
   U12571 : NOR2_X2 port map( A1 => n16527, A2 => n16534, ZN => n15916);
   U12572 : NOR2_X2 port map( A1 => n17411, A2 => n15588, ZN => n17677);
   U12573 : NOR2_X2 port map( A1 => n17074, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_3_port, ZN 
                           => pipeline_stageE_EXE_ALU_alu_shift_C86_n1);
   U12574 : AND2_X2 port map( A1 => pipeline_WB_controls_in_MEMWB_0_port, A2 =>
                           n17705, ZN => n14135);
   U12575 : XNOR2_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_add_29_n138, B 
                           => pipeline_stageD_evaluate_jump_target_add_29_n139,
                           ZN => pipeline_stageD_evaluate_jump_target_N38);
   U12576 : XNOR2_X1 port map( A => n17163, B => 
                           pipeline_stageD_evaluate_jump_target_add_29_n201, ZN
                           => pipeline_stageD_evaluate_jump_target_N47);
   U12577 : XNOR2_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_add_29_n191, B 
                           => n17169, ZN => 
                           pipeline_stageD_evaluate_jump_target_N50);
   U12578 : XNOR2_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_add_29_n172, B 
                           => pipeline_stageD_evaluate_jump_target_add_29_n175,
                           ZN => pipeline_stageD_evaluate_jump_target_N55);
   U12579 : XNOR2_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_add_29_n171, B 
                           => n17166, ZN => 
                           pipeline_stageD_evaluate_jump_target_N56);
   U12580 : XNOR2_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_add_29_n197, B 
                           => pipeline_stageD_evaluate_jump_target_add_29_n196,
                           ZN => pipeline_stageD_evaluate_jump_target_N48);
   U12581 : XNOR2_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_add_29_n144, B 
                           => n17182, ZN => 
                           pipeline_stageD_evaluate_jump_target_N36);
   U12582 : XNOR2_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_add_29_n165, B 
                           => n17164, ZN => 
                           pipeline_stageD_evaluate_jump_target_N58);
   U12583 : XNOR2_X1 port map( A => n17171, B => 
                           pipeline_stageD_evaluate_jump_target_add_29_n181, ZN
                           => pipeline_stageD_evaluate_jump_target_N53);
   U12584 : XNOR2_X1 port map( A => n17162, B => 
                           pipeline_stageD_evaluate_jump_target_add_29_n195, ZN
                           => pipeline_stageD_evaluate_jump_target_N49);
   U12585 : XNOR2_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_add_29_n177, B 
                           => n17179, ZN => 
                           pipeline_stageD_evaluate_jump_target_N54);
   U12586 : XNOR2_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_add_29_n126, B 
                           => n17175, ZN => 
                           pipeline_stageD_evaluate_jump_target_N42);
   U12587 : XNOR2_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_add_29_n132, B 
                           => pipeline_stageD_evaluate_jump_target_add_29_n133,
                           ZN => pipeline_stageD_evaluate_jump_target_N40);
   U12588 : XNOR2_X1 port map( A => n17161, B => 
                           pipeline_stageD_evaluate_jump_target_add_29_n150, ZN
                           => pipeline_stageD_evaluate_jump_target_N35);
   U12589 : XNOR2_X1 port map( A => n17168, B => 
                           pipeline_stageD_evaluate_jump_target_add_29_n189, ZN
                           => pipeline_stageD_evaluate_jump_target_N51);
   U12590 : XNOR2_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_add_29_n134, B 
                           => pipeline_stageD_evaluate_jump_target_add_29_n135,
                           ZN => pipeline_stageD_evaluate_jump_target_N39);
   U12591 : XNOR2_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_add_29_n160, B 
                           => pipeline_stageD_evaluate_jump_target_add_29_n163,
                           ZN => pipeline_stageD_evaluate_jump_target_N59);
   U12592 : XNOR2_X1 port map( A => n17173, B => 
                           pipeline_stageD_evaluate_jump_target_add_29_n213, ZN
                           => pipeline_stageD_evaluate_jump_target_N43);
   U12593 : XNOR2_X1 port map( A => n17165, B => 
                           pipeline_stageD_evaluate_jump_target_add_29_n169, ZN
                           => pipeline_stageD_evaluate_jump_target_N57);
   U12594 : NAND2_X1 port map( A1 => net175543, A2 => 
                           pipeline_nextPC_IFID_DEC_0_port, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n183);
   U12595 : AOI222_X1 port map( A1 => pipeline_nextPC_IFID_DEC_13_port, A2 => 
                           pipeline_stageD_offset_to_jump_temp_13_port, B1 => 
                           pipeline_nextPC_IFID_DEC_13_port, B2 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n202, C1
                           => pipeline_stageD_offset_to_jump_temp_13_port, C2 
                           => pipeline_stageD_evaluate_jump_target_add_29_n202,
                           ZN => n17163);
   U12596 : XNOR2_X1 port map( A => n17180, B => 
                           pipeline_stageD_evaluate_jump_target_add_29_n141, ZN
                           => pipeline_stageD_evaluate_jump_target_N37);
   U12597 : AOI22_X1 port map( A1 => pipeline_nextPC_IFID_DEC_2_port, A2 => 
                           pipeline_stageD_offset_to_jump_temp_2_port, B1 => 
                           n17404, B2 => n17470, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n150);
   U12598 : AOI222_X1 port map( A1 => pipeline_nextPC_IFID_DEC_23_port, A2 => 
                           pipeline_stageD_offset_to_jump_temp_23_port, B1 => 
                           pipeline_nextPC_IFID_DEC_23_port, B2 => n17166, C1 
                           => pipeline_stageD_offset_to_jump_temp_23_port, C2 
                           => n17166, ZN => n17165);
   U12599 : AOI222_X1 port map( A1 => pipeline_nextPC_IFID_DEC_17_port, A2 => 
                           pipeline_stageD_offset_to_jump_temp_17_port, B1 => 
                           pipeline_nextPC_IFID_DEC_17_port, B2 => n17169, C1 
                           => pipeline_stageD_evaluate_jump_target_add_29_n190,
                           C2 => pipeline_stageD_offset_to_jump_temp_17_port, 
                           ZN => n17168);
   U12600 : XNOR2_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_add_29_n185, B 
                           => pipeline_stageD_evaluate_jump_target_add_29_n182,
                           ZN => pipeline_stageD_evaluate_jump_target_N52);
   U12601 : AOI222_X1 port map( A1 => pipeline_nextPC_IFID_DEC_19_port, A2 => 
                           pipeline_stageD_offset_to_jump_temp_19_port, B1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n182, B2
                           => pipeline_nextPC_IFID_DEC_19_port, C1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n182, C2
                           => pipeline_stageD_offset_to_jump_temp_19_port, ZN 
                           => n17172);
   U12602 : AOI222_X1 port map( A1 => pipeline_nextPC_IFID_DEC_19_port, A2 => 
                           pipeline_stageD_offset_to_jump_temp_19_port, B1 => 
                           pipeline_nextPC_IFID_DEC_19_port, B2 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n182, C1
                           => pipeline_stageD_evaluate_jump_target_add_29_n182,
                           C2 => pipeline_stageD_offset_to_jump_temp_19_port, 
                           ZN => n17171);
   U12603 : AOI222_X1 port map( A1 => 
                           pipeline_stageD_offset_to_jump_temp_9_port, A2 => 
                           pipeline_nextPC_IFID_DEC_9_port, B1 => 
                           pipeline_stageD_offset_to_jump_temp_9_port, B2 => 
                           n17175, C1 => pipeline_nextPC_IFID_DEC_9_port, C2 =>
                           n17175, ZN => n17173);
   U12604 : XNOR2_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_add_29_n128, B 
                           => pipeline_stageD_evaluate_jump_target_add_29_n129,
                           ZN => pipeline_stageD_evaluate_jump_target_N41);
   U12605 : AOI222_X1 port map( A1 => pipeline_nextPC_IFID_DEC_11_port, A2 => 
                           pipeline_stageD_offset_to_jump_temp_11_port, B1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n208, B2
                           => pipeline_nextPC_IFID_DEC_11_port, C1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n208, C2
                           => pipeline_stageD_offset_to_jump_temp_11_port, ZN 
                           => n17178);
   U12606 : XNOR2_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_add_29_n203, B 
                           => pipeline_stageD_evaluate_jump_target_add_29_n202,
                           ZN => pipeline_stageD_evaluate_jump_target_N46);
   U12607 : AOI222_X1 port map( A1 => pipeline_nextPC_IFID_DEC_3_port, A2 => 
                           pipeline_stageD_offset_to_jump_temp_3_port, B1 => 
                           pipeline_nextPC_IFID_DEC_3_port, B2 => n17182, C1 =>
                           pipeline_stageD_offset_to_jump_temp_3_port, C2 => 
                           n17182, ZN => n17180);
   U12608 : AOI222_X1 port map( A1 => n17161, A2 => n17470, B1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n149, B2
                           => n17404, C1 => n17470, C2 => n17404, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n145);
   U12609 : NAND3_X1 port map( A1 => n17186, A2 => n17185, A3 => n17184, ZN => 
                           n17188);
   U12610 : XNOR2_X1 port map( A => n17192, B => n17191, ZN => 
                           pipeline_stageD_evaluate_jump_target_N62);
   U12611 : NAND2_X1 port map( A1 => n17190, A2 => n17189, ZN => n17192);
   U12612 : AOI21_X1 port map( B1 => n17201, B2 => n17451, A => n17200, ZN => 
                           n17202);
   U12613 : NAND2_X1 port map( A1 => n17166, A2 => 
                           pipeline_stageD_offset_to_jump_temp_23_port, ZN => 
                           n17195);
   U12614 : NAND2_X1 port map( A1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n170, A2
                           => pipeline_stageD_offset_to_jump_temp_23_port, ZN 
                           => n17194);
   U12615 : NAND3_X1 port map( A1 => n17196, A2 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n168, A3
                           => n17194, ZN => n17199);
   U12616 : NAND3_X1 port map( A1 => n17196, A2 => n17465, A3 => n17195, ZN => 
                           n17198);
   U12617 : NAND3_X1 port map( A1 => n17198, A2 => n17199, A3 => n17197, ZN => 
                           n17201);
   U12618 : NAND2_X1 port map( A1 => n17208, A2 => n17465, ZN => n17207);
   U12619 : NAND2_X1 port map( A1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n168, A2
                           => n17208, ZN => n17209);
   U12620 : OAI21_X1 port map( B1 => n17464, B2 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n174, A 
                           => pipeline_stageD_evaluate_jump_target_add_29_n172,
                           ZN => n17214);
   U12621 : AOI21_X1 port map( B1 => n17219, B2 => n17448, A => n17218, ZN => 
                           n17220);
   U12622 : NAND2_X1 port map( A1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n178, A2
                           => pipeline_stageD_evaluate_jump_target_add_29_n180,
                           ZN => n17217);
   U12623 : NAND2_X1 port map( A1 => n17172, A2 => n17463, ZN => n17216);
   U12624 : NAND3_X1 port map( A1 => n17216, A2 => n17217, A3 => n17215, ZN => 
                           n17219);
   U12625 : AOI222_X1 port map( A1 => pipeline_nextPC_IFID_DEC_19_port, A2 => 
                           pipeline_stageD_offset_to_jump_temp_19_port, B1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n182, B2
                           => pipeline_nextPC_IFID_DEC_19_port, C1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n182, C2
                           => pipeline_stageD_offset_to_jump_temp_19_port, ZN 
                           => pipeline_stageD_evaluate_jump_target_add_29_n178)
                           ;
   U12626 : NAND2_X1 port map( A1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n190, A2
                           => pipeline_stageD_offset_to_jump_temp_17_port, ZN 
                           => n17222);
   U12627 : OAI211_X1 port map( C1 => n17294, C2 => n17290, A => n17223, B => 
                           n17222, ZN => n17225);
   U12628 : NAND2_X1 port map( A1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n190, A2
                           => pipeline_nextPC_IFID_DEC_17_port, ZN => n17223);
   U12629 : OAI21_X1 port map( B1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n174, B2
                           => n17464, A => 
                           pipeline_stageD_evaluate_jump_target_add_29_n172, ZN
                           => n17227);
   U12630 : NAND2_X1 port map( A1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n196, A2
                           => pipeline_stageD_offset_to_jump_temp_15_port, ZN 
                           => n17230);
   U12631 : OAI21_X1 port map( B1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n196, B2
                           => pipeline_stageD_offset_to_jump_temp_15_port, A =>
                           pipeline_nextPC_IFID_DEC_15_port, ZN => n17231);
   U12632 : NAND2_X1 port map( A1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n196, A2
                           => pipeline_stageD_offset_to_jump_temp_15_port, ZN 
                           => n17232);
   U12633 : OAI21_X1 port map( B1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n196, B2
                           => pipeline_stageD_offset_to_jump_temp_15_port, A =>
                           pipeline_nextPC_IFID_DEC_15_port, ZN => n17233);
   U12634 : NAND2_X1 port map( A1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n178, A2
                           => pipeline_stageD_evaluate_jump_target_add_29_n180,
                           ZN => n17236);
   U12635 : NAND2_X1 port map( A1 => n17172, A2 => n17463, ZN => n17235);
   U12636 : NAND2_X1 port map( A1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n202, A2
                           => pipeline_stageD_offset_to_jump_temp_13_port, ZN 
                           => n17238);
   U12637 : OAI211_X1 port map( C1 => n17292, C2 => n17288, A => n17238, B => 
                           n17239, ZN => n17241);
   U12638 : NAND2_X1 port map( A1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n202, A2
                           => pipeline_nextPC_IFID_DEC_13_port, ZN => n17239);
   U12639 : NAND2_X1 port map( A1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n208, A2
                           => pipeline_stageD_offset_to_jump_temp_11_port, ZN 
                           => n17243);
   U12640 : OAI211_X1 port map( C1 => n17293, C2 => n17289, A => n17243, B => 
                           n17244, ZN => n17246);
   U12641 : NAND2_X1 port map( A1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n208, A2
                           => pipeline_nextPC_IFID_DEC_11_port, ZN => n17244);
   U12642 : OAI21_X1 port map( B1 => n17457, B2 => n17428, A => 
                           pipeline_stageD_evaluate_jump_target_add_29_n128, ZN
                           => n17251);
   U12643 : OAI22_X1 port map( A1 => n17255, A2 => n17254, B1 => 
                           pipeline_nextPC_IFID_DEC_10_port, B2 => 
                           pipeline_stageD_offset_to_jump_temp_10_port, ZN => 
                           n17256);
   U12644 : NAND2_X1 port map( A1 => n17176, A2 => 
                           pipeline_nextPC_IFID_DEC_9_port, ZN => n17248);
   U12645 : AOI21_X1 port map( B1 => n17176, B2 => 
                           pipeline_stageD_offset_to_jump_temp_9_port, A => 
                           n17247, ZN => n17249);
   U12646 : NAND3_X1 port map( A1 => n17251, A2 => 
                           pipeline_nextPC_IFID_DEC_9_port, A3 => n17250, ZN =>
                           n17253);
   U12647 : NAND3_X1 port map( A1 => n17253, A2 => n17440, A3 => n17252, ZN => 
                           n17254);
   U12648 : OAI21_X1 port map( B1 => n17428, B2 => n17457, A => 
                           pipeline_stageD_evaluate_jump_target_add_29_n128, ZN
                           => n17259);
   U12649 : NAND2_X1 port map( A1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n133, A2
                           => pipeline_stageD_offset_to_jump_temp_7_port, ZN =>
                           n17260);
   U12650 : OAI21_X1 port map( B1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n133, B2
                           => pipeline_stageD_offset_to_jump_temp_7_port, A => 
                           pipeline_nextPC_IFID_DEC_7_port, ZN => n17261);
   U12651 : OAI21_X1 port map( B1 => n17361, B2 => n17456, A => 
                           pipeline_stageD_evaluate_jump_target_add_29_n134, ZN
                           => n17263);
   U12652 : NAND2_X1 port map( A1 => pipeline_nextPC_IFID_DEC_5_port, A2 => 
                           pipeline_stageD_offset_to_jump_temp_5_port, ZN => 
                           n17266);
   U12653 : NAND2_X1 port map( A1 => pipeline_nextPC_IFID_DEC_5_port, A2 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n139, ZN
                           => n17265);
   U12654 : NAND2_X1 port map( A1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n139, A2
                           => pipeline_stageD_offset_to_jump_temp_5_port, ZN =>
                           n17264);
   U12655 : NAND2_X1 port map( A1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n145, A2
                           => pipeline_stageD_offset_to_jump_temp_3_port, ZN =>
                           n17269);
   U12656 : AOI21_X1 port map( B1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n145, B2
                           => pipeline_nextPC_IFID_DEC_3_port, A => n17291, ZN 
                           => n17270);
   U12657 : NAND2_X1 port map( A1 => n17181, A2 => 
                           pipeline_stageD_offset_to_jump_temp_3_port, ZN => 
                           n17267);
   U12658 : AOI21_X1 port map( B1 => n17181, B2 => 
                           pipeline_nextPC_IFID_DEC_3_port, A => n17291, ZN => 
                           n17268);
   U12659 : NAND3_X1 port map( A1 => n17268, A2 => n17455, A3 => n17267, ZN => 
                           n17273);
   U12660 : NAND3_X1 port map( A1 => n17270, A2 => n17412, A3 => n17269, ZN => 
                           n17271);
   U12661 : AOI222_X1 port map( A1 => pipeline_nextPC_IFID_DEC_1_port, A2 => 
                           pipeline_stageD_offset_to_jump_temp_1_port, B1 => 
                           n17167, B2 => pipeline_nextPC_IFID_DEC_1_port, C1 =>
                           pipeline_stageD_evaluate_jump_target_add_29_n214, C2
                           => pipeline_stageD_offset_to_jump_temp_1_port, ZN =>
                           n17274);
   U12662 : NAND2_X1 port map( A1 => net175543, A2 => 
                           pipeline_nextPC_IFID_DEC_0_port, ZN => n17275);
   U12663 : AOI21_X1 port map( B1 => n17406, B2 => n17275, A => n17446, ZN => 
                           n17277);
   U12664 : XNOR2_X1 port map( A => n17188, B => n17187, ZN => 
                           pipeline_stageD_evaluate_jump_target_N63);
   U12665 : NAND3_X1 port map( A1 => n17278, A2 => n17279, A3 => n17287, ZN => 
                           n17185);
   U12666 : NAND2_X1 port map( A1 => n17281, A2 => n17200, ZN => n17278);
   U12667 : NAND2_X1 port map( A1 => n17280, A2 => n17286, ZN => n17190);
   U12668 : XNOR2_X1 port map( A => n17280, B => 
                           pipeline_stageD_evaluate_jump_target_add_29_n157, ZN
                           => pipeline_stageD_evaluate_jump_target_N61);
   U12669 : NAND2_X1 port map( A1 => n17281, A2 => n17467, ZN => n17279);
   U12670 : NAND2_X1 port map( A1 => n17283, A2 => 
                           pipeline_stageD_offset_to_jump_temp_30_port, ZN => 
                           n17193);
   U12671 : XNOR2_X1 port map( A => n17283, B => 
                           pipeline_stageD_evaluate_jump_target_add_29_n159, ZN
                           => pipeline_stageD_evaluate_jump_target_N60);
   U12672 : OAI21_X1 port map( B1 => n17283, B2 => 
                           pipeline_stageD_offset_to_jump_temp_30_port, A => 
                           pipeline_nextPC_IFID_DEC_27_port, ZN => n17282);
   U12673 : NAND2_X1 port map( A1 => 
                           pipeline_stageD_offset_to_jump_temp_17_port, A2 => 
                           pipeline_nextPC_IFID_DEC_17_port, ZN => n17221);
   U12674 : NAND2_X1 port map( A1 => 
                           pipeline_stageD_offset_to_jump_temp_13_port, A2 => 
                           pipeline_nextPC_IFID_DEC_13_port, ZN => n17237);
   U12675 : NAND2_X1 port map( A1 => 
                           pipeline_stageD_offset_to_jump_temp_11_port, A2 => 
                           pipeline_nextPC_IFID_DEC_11_port, ZN => n17242);
   U12676 : NAND2_X1 port map( A1 => n17412, A2 => n17455, ZN => n17272);
   U12677 : NAND2_X1 port map( A1 => n17361, A2 => n17456, ZN => n17262);
   U12678 : NAND2_X1 port map( A1 => n17428, A2 => n17457, ZN => n17258);
   U12679 : NAND2_X1 port map( A1 => pipeline_stageD_offset_to_jump_temp_9_port
                           , A2 => pipeline_nextPC_IFID_DEC_9_port, ZN => 
                           n17252);
   U12680 : NAND2_X1 port map( A1 => n17458, A2 => n17252, ZN => n17247);
   U12681 : NAND2_X1 port map( A1 => n17428, A2 => n17457, ZN => n17250);
   U12682 : NAND2_X1 port map( A1 => n17444, A2 => n17459, ZN => n17245);
   U12683 : NAND2_X1 port map( A1 => n17445, A2 => n17460, ZN => n17240);
   U12684 : NAND2_X1 port map( A1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n188, A2
                           => n17462, ZN => n17224);
   U12685 : NAND2_X1 port map( A1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n180, A2
                           => n17463, ZN => n17234);
   U12686 : NAND2_X1 port map( A1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n180, A2
                           => n17463, ZN => n17215);
   U12687 : NAND2_X1 port map( A1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n174, A2
                           => n17464, ZN => n17213);
   U12688 : NAND2_X1 port map( A1 => 
                           pipeline_stageD_offset_to_jump_temp_23_port, A2 => 
                           pipeline_nextPC_IFID_DEC_23_port, ZN => n17208);
   U12689 : NAND2_X1 port map( A1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n174, A2
                           => n17464, ZN => n17226);
   U12690 : NAND2_X1 port map( A1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n168, A2
                           => n17465, ZN => n17210);
   U12691 : NAND2_X1 port map( A1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n168, A2
                           => n17465, ZN => n17197);
   U12692 : NAND2_X1 port map( A1 => n17200, A2 => n17467, ZN => n17183);
   U12693 : NAND2_X1 port map( A1 => 
                           pipeline_stageD_offset_to_jump_temp_30_port, A2 => 
                           pipeline_nextPC_IFID_DEC_29_port, ZN => n17184);
   U12694 : XNOR2_X1 port map( A => pipeline_stageD_offset_to_jump_temp_30_port
                           , B => pipeline_nextPC_IFID_DEC_30_port, ZN => 
                           n17187);
   U12695 : NAND2_X1 port map( A1 => n17200, A2 => n17467, ZN => n17189);
   U12696 : XNOR2_X1 port map( A => pipeline_stageD_offset_to_jump_temp_30_port
                           , B => n17452, ZN => n17191);
   U12697 : INV_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_add_29_n190, ZN
                           => n17170);
   U12698 : AND2_X1 port map( A1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n188, A2
                           => n17221, ZN => n17294);
   U12699 : AND2_X1 port map( A1 => n17221, A2 => n17462, ZN => n17290);
   U12700 : AND2_X1 port map( A1 => n17445, A2 => n17237, ZN => n17292);
   U12701 : AND2_X1 port map( A1 => n17460, A2 => n17237, ZN => n17288);
   U12702 : AND2_X1 port map( A1 => n17444, A2 => n17242, ZN => n17293);
   U12703 : AND2_X1 port map( A1 => n17459, A2 => n17242, ZN => n17289);
   U12704 : AND2_X1 port map( A1 => net175543, A2 => 
                           pipeline_nextPC_IFID_DEC_0_port, ZN => n17167);
   U12705 : AND2_X1 port map( A1 => net175543, A2 => 
                           pipeline_nextPC_IFID_DEC_0_port, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n214);
   U12706 : NOR2_X1 port map( A1 => n17406, A2 => n17275, ZN => n17276);
   U12707 : NOR2_X1 port map( A1 => n17277, A2 => n17276, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n149);
   U12708 : AND2_X1 port map( A1 => pipeline_stageD_offset_to_jump_temp_3_port,
                           A2 => pipeline_nextPC_IFID_DEC_3_port, ZN => n17291)
                           ;
   U12709 : AND3_X1 port map( A1 => n17266, A2 => n17265, A3 => n17264, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n134);
   U12710 : AND2_X1 port map( A1 => n17259, A2 => n17258, ZN => n17176);
   U12711 : AND2_X1 port map( A1 => n17249, A2 => n17248, ZN => n17257);
   U12712 : AND2_X1 port map( A1 => n17177, A2 => 
                           pipeline_stageD_offset_to_jump_temp_9_port, ZN => 
                           n17255);
   U12713 : AND3_X1 port map( A1 => n17231, A2 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n194, A3
                           => n17230, ZN => n17229);
   U12714 : AND2_X1 port map( A1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n194, A2
                           => n17461, ZN => n17228);
   U12715 : AND3_X1 port map( A1 => n17236, A2 => n17235, A3 => n17234, ZN => 
                           n17179);
   U12716 : INV_X1 port map( A => pipeline_stageD_offset_to_jump_temp_21_port, 
                           ZN => n17218);
   U12717 : AND2_X1 port map( A1 => n17166, A2 => 
                           pipeline_stageD_offset_to_jump_temp_23_port, ZN => 
                           n17203);
   U12718 : AND2_X1 port map( A1 => n17166, A2 => 
                           pipeline_nextPC_IFID_DEC_23_port, ZN => n17204);
   U12719 : OR3_X1 port map( A1 => n17203, A2 => n17204, A3 => n17207, ZN => 
                           n17212);
   U12720 : AND2_X1 port map( A1 => n17227, A2 => n17226, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n170);
   U12721 : AND2_X1 port map( A1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n170, A2
                           => pipeline_nextPC_IFID_DEC_23_port, ZN => n17205);
   U12722 : AND2_X1 port map( A1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n170, A2
                           => pipeline_stageD_offset_to_jump_temp_23_port, ZN 
                           => n17206);
   U12723 : OR3_X1 port map( A1 => n17205, A2 => n17206, A3 => n17209, ZN => 
                           n17211);
   U12724 : AND3_X1 port map( A1 => n17212, A2 => n17211, A3 => n17210, ZN => 
                           n17164);
   U12725 : INV_X1 port map( A => pipeline_stageD_offset_to_jump_temp_30_port, 
                           ZN => n17200);
   U12726 : OR2_X1 port map( A1 => n17200, A2 => n17466, ZN => n17285);
   U12727 : AND2_X1 port map( A1 => n17200, A2 => n17466, ZN => n17284);
   U12728 : AND2_X1 port map( A1 => n17282, A2 => n17193, ZN => n17281);
   U12729 : AND2_X1 port map( A1 => n17183, A2 => 
                           pipeline_stageD_offset_to_jump_temp_30_port, ZN => 
                           n17287);
   U12730 : AND2_X1 port map( A1 => n17282, A2 => n17193, ZN => n17280);
   U12731 : OR2_X1 port map( A1 => n17200, A2 => n17467, ZN => n17286);
   U12732 : INV_X1 port map( A => n17170, ZN => n17169);
   U12733 : CLKBUF_X1 port map( A => 
                           pipeline_stageD_evaluate_jump_target_add_29_n208, Z 
                           => n17174);
   U12734 : CLKBUF_X1 port map( A => n17177, Z => n17175);
   U12735 : CLKBUF_X1 port map( A => n17181, Z => n17182);
   U12736 : AOI222_X2 port map( A1 => n17274, A2 => n17470, B1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n149, B2
                           => n17404, C1 => n17470, C2 => n17404, ZN => n17181)
                           ;
   U12737 : NOR2_X2 port map( A1 => n17257, A2 => n17256, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n208);
   U12738 : AND2_X2 port map( A1 => n17225, A2 => n17224, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n182);
   U12739 : AND2_X2 port map( A1 => n17214, A2 => n17213, ZN => n17166);
   U12740 : AND2_X2 port map( A1 => n17241, A2 => n17240, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n196);
   U12741 : AOI21_X1 port map( B1 => 
                           pipeline_stageD_evaluate_jump_target_add_29_n160, B2
                           => n17285, A => n17284, ZN => n17283);
   U12742 : AND2_X2 port map( A1 => n17246, A2 => n17245, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n202);
   U12743 : AND3_X2 port map( A1 => n17273, A2 => n17272, A3 => n17271, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n139);
   U12744 : AOI21_X2 port map( B1 => n17179, B2 => 
                           pipeline_nextPC_IFID_DEC_21_port, A => n17220, ZN =>
                           pipeline_stageD_evaluate_jump_target_add_29_n172);
   U12745 : AOI211_X2 port map( C1 => n17162, C2 => n17461, A => n17229, B => 
                           n17228, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n190);
   U12746 : AND2_X2 port map( A1 => n17261, A2 => n17260, ZN => 
                           pipeline_stageD_evaluate_jump_target_add_29_n128);
   U12747 : OR2_X1 port map( A1 => n17428, A2 => n17457, ZN => n17295);
   U12748 : AND2_X1 port map( A1 => pipeline_stageE_EXE_ALU_alu_shift_N202, A2 
                           => n17742, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C88_ML_int_1_0_port);
   U12749 : NAND2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_1_port, A2 
                           => n17742, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n46);
   U12750 : NOR2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, A2 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_SH_1_port, 
                           ZN => pipeline_stageE_EXE_ALU_alu_shift_C50_n50);
   U12751 : NOR2_X1 port map( A1 => n17742, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_1_port, ZN 
                           => pipeline_stageE_EXE_ALU_alu_shift_C50_n49);
   U12752 : NOR2_X1 port map( A1 => n17739, A2 => n17074, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n76);
   U12753 : AOI22_X1 port map( A1 => pipeline_stageE_input1_to_ALU_1_port, A2 
                           => pipeline_stageE_EXE_ALU_alu_shift_C86_n26, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N202, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n27, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n151);
   U12754 : NOR2_X1 port map( A1 => n17081, A2 => n17296, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n73);
   U12755 : INV_X1 port map( A => pipeline_stageE_EXE_ALU_alu_shift_C50_n46, ZN
                           => pipeline_stageE_EXE_ALU_alu_shift_C50_n167);
   U12756 : INV_X1 port map( A => n17739, ZN => n17296);
   U12757 : INV_X1 port map( A => n17112, ZN => n17297);
   U12758 : INV_X1 port map( A => pipeline_stageE_EXE_ALU_alu_shift_C50_n124, 
                           ZN => pipeline_stageE_EXE_ALU_alu_shift_C50_n72);
   U12759 : AND2_X1 port map( A1 => n17074, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n148, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n10);
   U12760 : AND2_X1 port map( A1 => pipeline_stageE_EXE_ALU_alu_shift_C50_n148,
                           A2 => n17081, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C50_n8);
   U12761 : NOR2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, A2 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_SH_1_port, 
                           ZN => pipeline_stageE_EXE_ALU_alu_shift_C86_n27);
   U12762 : NOR2_X1 port map( A1 => n17742, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_1_port, ZN 
                           => pipeline_stageE_EXE_ALU_alu_shift_C86_n26);
   U12763 : AOI222_X1 port map( A1 => n17111, A2 => n12649, B1 => 
                           pipeline_stageE_input1_to_ALU_1_port, B2 => n17110, 
                           C1 => pipeline_stageE_EXE_ALU_alu_shift_N202, C2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_1_port, ZN 
                           => pipeline_stageE_EXE_ALU_alu_shift_C86_n170);
   U12764 : NAND2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_3_port, A2 
                           => pipeline_stageE_EXE_ALU_alu_shift_N202, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n104);
   U12765 : NAND2_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, A2 
                           => pipeline_stageE_EXE_ALU_alu_shift_N202, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n4);
   U12766 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port, ZN 
                           => n17302);
   U12767 : AND2_X1 port map( A1 => n17074, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_3_port, ZN 
                           => pipeline_stageE_EXE_ALU_alu_shift_C86_n136);
   U12768 : AND2_X1 port map( A1 => pipeline_stageE_EXE_ALU_alu_shift_C86_n131,
                           A2 => n17074, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n15);
   U12769 : AND2_X1 port map( A1 => pipeline_stageE_EXE_ALU_alu_shift_C86_n131,
                           A2 => n17081, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C86_n19);
   U12770 : AOI22_X1 port map( A1 => pipeline_stageE_input1_to_ALU_1_port, A2 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_n51, B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N202, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n52, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n160);
   U12771 : INV_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_1_port, ZN 
                           => n17303);
   U12772 : NOR2_X1 port map( A1 => n17303, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, ZN 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_n2);
   U12773 : AND2_X1 port map( A1 => n17074, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_3_port, ZN 
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_n105);
   U12774 : AND2_X1 port map( A1 => n17074, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n158, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n12);
   U12775 : AND2_X1 port map( A1 => pipeline_stageE_EXE_ALU_alu_shift_C48_n158,
                           A2 => n17081, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_n10);
   U12776 : OAI21_X1 port map( B1 => n15218, B2 => n15220, A => n15221, ZN => 
                           n15205);
   U12777 : INV_X4 port map( A => n17737, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_4_port);
   U12778 : CLKBUF_X1 port map( A => n13172, Z => n17706);
   U12779 : CLKBUF_X1 port map( A => n13166, Z => n17708);
   U12780 : CLKBUF_X1 port map( A => n13160, Z => n17710);
   U12781 : CLKBUF_X1 port map( A => n13154, Z => n17712);
   U12782 : CLKBUF_X1 port map( A => n13148, Z => n17714);
   U12783 : CLKBUF_X1 port map( A => n13142, Z => n17716);
   U12784 : CLKBUF_X1 port map( A => n13136, Z => n17718);
   U12785 : CLKBUF_X1 port map( A => n13130, Z => n17720);
   U12786 : CLKBUF_X1 port map( A => n13124, Z => n17722);
   U12787 : CLKBUF_X1 port map( A => n13118, Z => n17724);
   U12788 : CLKBUF_X1 port map( A => n13112, Z => n17726);
   U12789 : CLKBUF_X1 port map( A => n13106, Z => n17728);
   U12790 : CLKBUF_X1 port map( A => n13169, Z => n17707);
   U12791 : CLKBUF_X1 port map( A => n13163, Z => n17709);
   U12792 : CLKBUF_X1 port map( A => n13157, Z => n17711);
   U12793 : CLKBUF_X1 port map( A => n13145, Z => n17715);
   U12794 : CLKBUF_X1 port map( A => n13139, Z => n17717);
   U12795 : CLKBUF_X1 port map( A => n13133, Z => n17719);
   U12796 : CLKBUF_X1 port map( A => n13127, Z => n17721);
   U12797 : CLKBUF_X1 port map( A => n13121, Z => n17723);
   U12798 : CLKBUF_X1 port map( A => n13115, Z => n17725);
   U12799 : CLKBUF_X1 port map( A => n13109, Z => n17727);
   U12800 : CLKBUF_X1 port map( A => n13097, Z => n17731);
   U12801 : CLKBUF_X1 port map( A => n13082, Z => n17736);
   U12802 : CLKBUF_X1 port map( A => n13088, Z => n17734);
   U12803 : CLKBUF_X1 port map( A => n13094, Z => n17732);
   U12804 : CLKBUF_X1 port map( A => n13085, Z => n17735);
   U12805 : CLKBUF_X1 port map( A => n13100, Z => n17730);
   U12806 : CLKBUF_X1 port map( A => n13091, Z => n17733);
   U12807 : INV_X1 port map( A => n15116, ZN => n13184);
   U12808 : INV_X1 port map( A => n15120, ZN => n13178);
   U12809 : INV_X1 port map( A => n15104, ZN => n13202);
   U12810 : INV_X1 port map( A => n15112, ZN => n13190);
   U12811 : INV_X1 port map( A => n15114, ZN => n13187);
   U12812 : INV_X1 port map( A => n15102, ZN => n13205);
   U12813 : INV_X1 port map( A => n15108, ZN => n13196);
   U12814 : INV_X1 port map( A => n15110, ZN => n13193);
   U12815 : INV_X1 port map( A => n15118, ZN => n13181);
   U12816 : INV_X1 port map( A => n15084, ZN => n13232);
   U12817 : INV_X1 port map( A => n15122, ZN => n13175);
   U12818 : INV_X1 port map( A => n15096, ZN => n13214);
   U12819 : INV_X1 port map( A => n15092, ZN => n13220);
   U12820 : INV_X1 port map( A => n15088, ZN => n13226);
   U12821 : INV_X1 port map( A => n15106, ZN => n13199);
   U12822 : INV_X1 port map( A => n15064, ZN => n13262);
   U12823 : INV_X1 port map( A => n15080, ZN => n13238);
   U12824 : INV_X1 port map( A => n15094, ZN => n13217);
   U12825 : INV_X1 port map( A => n15076, ZN => n13244);
   U12826 : INV_X1 port map( A => n15090, ZN => n13223);
   U12827 : INV_X1 port map( A => n15072, ZN => n13250);
   U12828 : INV_X1 port map( A => n15082, ZN => n13235);
   U12829 : INV_X1 port map( A => n15068, ZN => n13256);
   U12830 : INV_X1 port map( A => n14988, ZN => n13268);
   U12831 : INV_X1 port map( A => n15062, ZN => n13265);
   U12832 : INV_X1 port map( A => n15100, ZN => n13208);
   U12833 : INV_X1 port map( A => n15086, ZN => n13229);
   U12834 : INV_X1 port map( A => n15074, ZN => n13247);
   U12835 : INV_X1 port map( A => n15098, ZN => n13211);
   U12836 : INV_X1 port map( A => n15078, ZN => n13241);
   U12837 : INV_X1 port map( A => n15066, ZN => n13259);
   U12838 : INV_X1 port map( A => n15070, ZN => n13253);
   U12839 : INV_X1 port map( A => n17420, ZN => n17682);
   U12840 : AND2_X1 port map( A1 => n14167, A2 => n14947, ZN => n17420);
   U12841 : AND2_X1 port map( A1 => pipeline_EXE_controls_in_IDEX_8_port, A2 =>
                           pipeline_IDEX_Stage_N181, ZN => 
                           pipeline_IDEX_Stage_N197);
   U12842 : INV_X1 port map( A => n15621, ZN => n3987);
   U12843 : AND3_X1 port map( A1 => n17625, A2 => n17626, A3 => n17627, ZN => 
                           n17635);
   U12844 : OR2_X1 port map( A1 => pipeline_stageE_EXE_ALU_alu_shift_N202, A2 
                           => pipeline_EXE_controls_in_EXEcute_4_port, ZN => 
                           n17633);
   U12845 : OR2_X1 port map( A1 => pipeline_stageE_EXE_ALU_alu_shift_N202, A2 
                           => pipeline_EXE_controls_in_EXEcute_3_port, ZN => 
                           n17634);
   U12846 : AND2_X1 port map( A1 => n14995, A2 => 
                           pipeline_EXE_controls_in_EXEcute_6_port, ZN => 
                           n17529);
   U12847 : INV_X1 port map( A => n15005, ZN => n15001);
   U12848 : AND2_X1 port map( A1 => n15165, A2 => n15166, ZN => n17540);
   U12849 : INV_X1 port map( A => n15007, ZN => n17551);
   U12850 : AND2_X1 port map( A1 => n15145, A2 => n15138, ZN => n17615);
   U12851 : AND3_X1 port map( A1 => n17546, A2 => n15009, A3 => n15010, ZN => 
                           n17547);
   U12852 : INV_X1 port map( A => n15161, ZN => n15138);
   U12853 : INV_X1 port map( A => n15164, ZN => n15165);
   U12854 : AND2_X1 port map( A1 => n15011, A2 => n17533, ZN => n17546);
   U12855 : AND2_X1 port map( A1 => n15597, A2 => n15049, ZN => n15058);
   U12856 : INV_X1 port map( A => n15445, ZN => n15429);
   U12857 : INV_X1 port map( A => n15268, ZN => n15281);
   U12858 : INV_X1 port map( A => n17649, ZN => n15335);
   U12859 : INV_X1 port map( A => n15282, ZN => n15267);
   U12860 : INV_X1 port map( A => n15015, ZN => n17535);
   U12861 : AND3_X1 port map( A1 => n17609, A2 => n17610, A3 => n17611, ZN => 
                           n17539);
   U12862 : AND2_X1 port map( A1 => pipeline_stageE_input1_to_ALU_25_port, A2 
                           => n15234, ZN => n17604);
   U12863 : AND2_X1 port map( A1 => n15235, A2 => n15234, ZN => n17605);
   U12864 : AND2_X1 port map( A1 => n15235, A2 => 
                           pipeline_stageE_input1_to_ALU_25_port, ZN => n17606)
                           ;
   U12865 : NAND2_X1 port map( A1 => n17593, A2 => n17594, ZN => n15282);
   U12866 : INV_X1 port map( A => n17598, ZN => n17596);
   U12867 : INV_X1 port map( A => n15314, ZN => n15332);
   U12868 : INV_X1 port map( A => n16631, ZN => n16630);
   U12869 : INV_X1 port map( A => n17738, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_A_16_port);
   U12870 : INV_X1 port map( A => pipeline_stageE_input1_to_ALU_16_port, ZN => 
                           n17738);
   U12871 : AND2_X1 port map( A1 => n17101, A2 => n15397, ZN => n17592);
   U12872 : OR2_X1 port map( A1 => n17101, A2 => n15397, ZN => n17591);
   U12873 : OR2_X1 port map( A1 => n15461, A2 => n15480, ZN => n17586);
   U12874 : INV_X1 port map( A => n15461, ZN => n17587);
   U12875 : NAND2_X1 port map( A1 => n15478, A2 => n15479, ZN => n15494);
   U12876 : OR2_X1 port map( A1 => pipeline_stageE_input1_to_ALU_7_port, A2 => 
                           n15521, ZN => n17583);
   U12877 : AND2_X1 port map( A1 => n15525, A2 => n15540, ZN => n17584);
   U12878 : AND3_X1 port map( A1 => n17568, A2 => n17569, A3 => n17570, ZN => 
                           pipeline_stageE_input2_to_ALU_0_port);
   U12879 : NOR2_X1 port map( A1 => n17387, A2 => n14982, ZN => n17665);
   U12880 : OR2_X1 port map( A1 => n17575, A2 => n17573, ZN => 
                           pipeline_stageE_EXE_ALU_alu_shift_N202);
   U12881 : AND2_X1 port map( A1 => n16620, A2 => n13965, ZN => n17575);
   U12882 : OR2_X1 port map( A1 => n16693, A2 => 
                           pipeline_stageE_input1_to_ALU_1_port, ZN => n15050);
   U12883 : AND2_X1 port map( A1 => n17740, A2 => n17381, ZN => n17576);
   U12884 : INV_X1 port map( A => n17641, ZN => n17642);
   U12885 : INV_X1 port map( A => n16619, ZN => n17572);
   U12886 : OR2_X1 port map( A1 => n16796, A2 => n16795, ZN => n17558);
   U12887 : INV_X1 port map( A => n16607, ZN => n17667);
   U12888 : AND2_X1 port map( A1 => pipeline_Reg2_Addr_to_exe_3_port, A2 => 
                           n17385, ZN => n17549);
   U12889 : AND2_X1 port map( A1 => n17314, A2 => 
                           pipeline_Reg2_Addr_to_exe_0_port, ZN => n17548);
   U12890 : INV_X1 port map( A => n17346, ZN => n17666);
   U12891 : OR2_X1 port map( A1 => n14982, A2 => n17387, ZN => n17346);
   U12892 : OR3_X1 port map( A1 => n16785, A2 => n16786, A3 => n16554, ZN => 
                           n14982);
   U12893 : INV_X1 port map( A => n17555, ZN => n17553);
   U12894 : AND3_X1 port map( A1 => n17637, A2 => n17638, A3 => n17639, ZN => 
                           n17402);
   U12895 : INV_X1 port map( A => n14885, ZN => n17640);
   U12896 : AND4_X1 port map( A1 => n17644, A2 => n17645, A3 => n17646, A4 => 
                           n17647, ZN => n16554);
   U12897 : AND2_X1 port map( A1 => n17340, A2 => n17393, ZN => n17647);
   U12898 : INV_X1 port map( A => n16585, ZN => n16561);
   U12899 : INV_X1 port map( A => n16586, ZN => n16805);
   U12900 : NOR2_X1 port map( A1 => n16666, A2 => 
                           pipeline_stageE_input1_to_ALU_10_port, ZN => n15461)
                           ;
   U12901 : NOR2_X1 port map( A1 => n14168, A2 => n15833, ZN => n15610);
   U12902 : NOR2_X1 port map( A1 => n15829, A2 => n15828, ZN => n17332);
   U12903 : NOR2_X1 port map( A1 => n15827, A2 => n15828, ZN => n17330);
   U12904 : NOR2_X1 port map( A1 => n15829, A2 => n15828, ZN => n17333);
   U12905 : NOR2_X1 port map( A1 => n15827, A2 => n15828, ZN => n17331);
   U12906 : OAI21_X1 port map( B1 => n17666, B2 => n17123, A => n17327, ZN => 
                           n16777);
   U12907 : NOR2_X1 port map( A1 => n14863, A2 => n14878, ZN => n14250);
   U12908 : NOR2_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_3_port, A2
                           => n15584, ZN => n14964);
   U12909 : NOR2_X1 port map( A1 => n16608, A2 => n17083, ZN => n15161);
   U12910 : NOR4_X1 port map( A1 => n16778, A2 => n16561, A3 => n16779, A4 => 
                           n16780, ZN => n17669);
   U12911 : NOR2_X1 port map( A1 => Rst, A2 => n15646, ZN => n15611);
   U12912 : OAI21_X1 port map( B1 => n16583, B2 => n16588, A => n17703, ZN => 
                           n13106);
   U12913 : OAI21_X1 port map( B1 => n16581, B2 => n16588, A => n17704, ZN => 
                           n13112);
   U12914 : OAI21_X1 port map( B1 => n16579, B2 => n16588, A => n17701, ZN => 
                           n13118);
   U12915 : OAI21_X1 port map( B1 => n16576, B2 => n16588, A => n17704, ZN => 
                           n13124);
   U12916 : OAI21_X1 port map( B1 => n16583, B2 => n16587, A => n17703, ZN => 
                           n13130);
   U12917 : OAI21_X1 port map( B1 => n16581, B2 => n16587, A => n17703, ZN => 
                           n13136);
   U12918 : OAI21_X1 port map( B1 => n16579, B2 => n16587, A => n17703, ZN => 
                           n13142);
   U12919 : OAI21_X1 port map( B1 => n16576, B2 => n16587, A => n17703, ZN => 
                           n13148);
   U12920 : OAI21_X1 port map( B1 => n16583, B2 => n16577, A => n17705, ZN => 
                           n13154);
   U12921 : OAI21_X1 port map( B1 => n16581, B2 => n16577, A => n17705, ZN => 
                           n13160);
   U12922 : OAI21_X1 port map( B1 => n16579, B2 => n16577, A => n17705, ZN => 
                           n13166);
   U12923 : OAI21_X1 port map( B1 => n16576, B2 => n16577, A => n17705, ZN => 
                           n13172);
   U12924 : OAI21_X1 port map( B1 => n16578, B2 => n16577, A => n17705, ZN => 
                           n13169);
   U12925 : OAI21_X1 port map( B1 => n16580, B2 => n16577, A => n17705, ZN => 
                           n13163);
   U12926 : OAI21_X1 port map( B1 => n16582, B2 => n16577, A => n17703, ZN => 
                           n13157);
   U12927 : NAND2_X1 port map( A1 => n16584, A2 => n17643, ZN => n16577);
   U12928 : OAI21_X1 port map( B1 => n16586, B2 => n16587, A => n17705, ZN => 
                           n13151);
   U12929 : OAI21_X1 port map( B1 => n16578, B2 => n16587, A => n17703, ZN => 
                           n13145);
   U12930 : OAI21_X1 port map( B1 => n16580, B2 => n16587, A => n17704, ZN => 
                           n13139);
   U12931 : OAI21_X1 port map( B1 => n16582, B2 => n16587, A => n17703, ZN => 
                           n13133);
   U12932 : OAI21_X1 port map( B1 => n16586, B2 => n16588, A => n17703, ZN => 
                           n13127);
   U12933 : OAI21_X1 port map( B1 => n16578, B2 => n16588, A => n17704, ZN => 
                           n13121);
   U12934 : OAI21_X1 port map( B1 => n16580, B2 => n16588, A => n17702, ZN => 
                           n13115);
   U12935 : OAI21_X1 port map( B1 => n16582, B2 => n16588, A => n17704, ZN => 
                           n13109);
   U12936 : OAI21_X1 port map( B1 => n16586, B2 => n16589, A => n17704, ZN => 
                           n13103);
   U12937 : OAI21_X1 port map( B1 => n16589, B2 => n16578, A => n17704, ZN => 
                           n13097);
   U12938 : NAND2_X1 port map( A1 => n17703, A2 => n17650, ZN => n13058);
   U12939 : OAI21_X1 port map( B1 => n16583, B2 => n16589, A => n17704, ZN => 
                           n13082);
   U12940 : OAI21_X1 port map( B1 => n16589, B2 => n16581, A => n17704, ZN => 
                           n13088);
   U12941 : NAND2_X1 port map( A1 => n17703, A2 => n17651, ZN => n13061);
   U12942 : NAND2_X1 port map( A1 => n17703, A2 => n17657, ZN => n13073);
   U12943 : NAND2_X1 port map( A1 => n17703, A2 => n17661, ZN => n13079);
   U12944 : OAI21_X1 port map( B1 => n16589, B2 => n16579, A => n17704, ZN => 
                           n13094);
   U12945 : OAI21_X1 port map( B1 => n16589, B2 => n16582, A => n17704, ZN => 
                           n13085);
   U12946 : NAND2_X1 port map( A1 => n17703, A2 => n17658, ZN => n13076);
   U12947 : NAND2_X1 port map( A1 => n17703, A2 => n17656, ZN => n13070);
   U12948 : OAI21_X1 port map( B1 => n16589, B2 => n16576, A => n17704, ZN => 
                           n13100);
   U12949 : NAND2_X1 port map( A1 => n17703, A2 => n17655, ZN => n13067);
   U12950 : OAI21_X1 port map( B1 => n16589, B2 => n16580, A => n17704, ZN => 
                           n13091);
   U12951 : NAND2_X1 port map( A1 => n17703, A2 => n17654, ZN => n13064);
   U12952 : NAND2_X1 port map( A1 => n16819, A2 => n17098, ZN => n16594);
   U12953 : NAND2_X1 port map( A1 => n16822, A2 => n17098, ZN => n16593);
   U12954 : NAND2_X1 port map( A1 => n16821, A2 => n17098, ZN => n16592);
   U12955 : NAND2_X1 port map( A1 => n17660, A2 => n17098, ZN => n16590);
   U12956 : NAND2_X1 port map( A1 => n16817, A2 => n17098, ZN => n16596);
   U12957 : NAND2_X1 port map( A1 => n17125, A2 => n17098, ZN => n16597);
   U12958 : NOR2_X1 port map( A1 => n14863, A2 => n14866, ZN => n14213);
   U12959 : NOR2_X1 port map( A1 => n14864, A2 => n14867, ZN => n14215);
   U12960 : NOR2_X1 port map( A1 => n14864, A2 => n14873, ZN => n14233);
   U12961 : NOR2_X1 port map( A1 => n14865, A2 => n14873, ZN => n14235);
   U12962 : NOR2_X1 port map( A1 => n14863, A2 => n14872, ZN => n14238);
   U12963 : NOR2_X1 port map( A1 => n14863, A2 => n14873, ZN => n14237);
   U12964 : NOR2_X1 port map( A1 => n14878, A2 => n14864, ZN => n14240);
   U12965 : NOR2_X1 port map( A1 => n14865, A2 => n14878, ZN => n14248);
   U12966 : NOR2_X1 port map( A1 => n14865, A2 => n14879, ZN => n14247);
   U12967 : NOR2_X1 port map( A1 => n14879, A2 => n14863, ZN => n14249);
   U12968 : NAND3_X1 port map( A1 => n17704, A2 => n17421, A3 => 
                           pipeline_EXE_controls_in_EXEcute_5_port, ZN => 
                           n14949);
   U12969 : INV_X2 port map( A => Rst, ZN => n17705);
   U12970 : NOR3_X1 port map( A1 => n15830, A2 => n15832, A3 => n15828, ZN => 
                           n15608);
   U12971 : AOI221_X1 port map( B1 => 
                           pipeline_stageD_offset_to_jump_temp_1_port, B2 => 
                           n14044, C1 => net175543, C2 => n14044, A => n14065, 
                           ZN => n14006);
   U12972 : NOR2_X1 port map( A1 => n14862, A2 => n14863, ZN => n17354);
   U12973 : NOR2_X1 port map( A1 => n14862, A2 => n14864, ZN => n17353);
   U12974 : NOR2_X1 port map( A1 => n14860, A2 => n14867, ZN => n17351);
   U12975 : NOR2_X1 port map( A1 => n14865, A2 => n14867, ZN => n17357);
   U12976 : NOR2_X1 port map( A1 => n14862, A2 => n14863, ZN => n17356);
   U12977 : NOR2_X1 port map( A1 => n14862, A2 => n14864, ZN => n17355);
   U12978 : NOR2_X1 port map( A1 => n14860, A2 => n14867, ZN => n17352);
   U12979 : NOR2_X1 port map( A1 => n14865, A2 => n14867, ZN => n17358);
   U12980 : NOR2_X1 port map( A1 => n14862, A2 => n14863, ZN => n17368);
   U12981 : NOR2_X1 port map( A1 => n14862, A2 => n14864, ZN => n17367);
   U12982 : AOI221_X1 port map( B1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_1_port, B2 
                           => n14968, C1 => n17741, C2 => n14981, A => n17103, 
                           ZN => n14975);
   U12983 : NOR2_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_2_port, A2
                           => n15581, ZN => n17359);
   U12984 : NAND2_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_4_port, 
                           A2 => n15573, ZN => n17678);
   U12985 : NOR2_X1 port map( A1 => n17405, A2 => n15581, ZN => n17360);
   U12986 : NAND2_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_4_port, 
                           A2 => n15573, ZN => n17679);
   U12987 : NOR2_X1 port map( A1 => n15834, A2 => n14127, ZN => n17676);
   U12988 : NAND2_X1 port map( A1 => n17674, A2 => n13944, ZN => n17622);
   U12989 : NAND2_X1 port map( A1 => pipeline_stageF_PC_plus4_N36, A2 => n17108
                           , ZN => n17621);
   U12990 : AOI21_X1 port map( B1 => n17631, B2 => n17632, A => 
                           pipeline_EXE_controls_in_EXEcute_6_port, ZN => 
                           n17630);
   U12991 : OAI211_X1 port map( C1 => n17119, C2 => 
                           pipeline_EXE_controls_in_EXEcute_2_port, A => n17742
                           , B => n17633, ZN => n17632);
   U12992 : OAI211_X1 port map( C1 => n17119, C2 => 
                           pipeline_stageE_EXE_ALU_add_alu_sCout_0_port, A => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, B 
                           => n17634, ZN => n17631);
   U12993 : NOR2_X1 port map( A1 => n17405, A2 => n15581, ZN => n17681);
   U12994 : NOR2_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_2_port, A2
                           => n15581, ZN => n17680);
   U12995 : AOI21_X1 port map( B1 => n15005, B2 => 
                           pipeline_EXE_controls_in_EXEcute_4_port, A => n17528
                           , ZN => n17618);
   U12996 : NOR2_X1 port map( A1 => n15161, A2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N136, ZN => n17608
                           );
   U12997 : XNOR2_X1 port map( A => n17104, B => n15137, ZN => n17614);
   U12998 : AOI21_X1 port map( B1 => n17617, B2 => n15142, A => n15161, ZN => 
                           n17616);
   U12999 : NAND2_X1 port map( A1 => n15146, A2 => n15147, ZN => n17617);
   U13000 : NAND2_X1 port map( A1 => n15165, A2 => n15147, ZN => n17612);
   U13001 : AOI221_X1 port map( B1 => pipeline_stageE_input1_to_ALU_19_port, B2
                           => n15314, C1 => n17649, C2 => n15316, A => n15317, 
                           ZN => n15296);
   U13002 : NAND2_X1 port map( A1 => pipeline_stageE_input1_to_ALU_27_port, A2 
                           => n15204, ZN => n17611);
   U13003 : NOR2_X1 port map( A1 => pipeline_stageE_input1_to_ALU_23_port, A2 
                           => n15263, ZN => n17603);
   U13004 : AOI21_X1 port map( B1 => n17595, B2 => n17596, A => n17597, ZN => 
                           n17594);
   U13005 : OAI21_X1 port map( B1 => n15301, B2 => n15297, A => n15299, ZN => 
                           n17597);
   U13006 : NAND2_X1 port map( A1 => n15319, A2 => n17599, ZN => n17595);
   U13007 : NAND2_X1 port map( A1 => n15314, A2 => 
                           pipeline_stageE_input1_to_ALU_19_port, ZN => n17599)
                           ;
   U13008 : NOR2_X1 port map( A1 => n17601, A2 => n17598, ZN => n17600);
   U13009 : NAND2_X1 port map( A1 => n15316, A2 => n17602, ZN => n17598);
   U13010 : NOR2_X1 port map( A1 => n15301, A2 => n15298, ZN => n17602);
   U13011 : NAND2_X1 port map( A1 => pipeline_stageE_input1_to_ALU_11_port, A2 
                           => n15459, ZN => n17590);
   U13012 : NAND2_X1 port map( A1 => pipeline_stageE_input1_to_ALU_7_port, A2 
                           => n15521, ZN => n17581);
   U13013 : NAND2_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_0_port, 
                           A2 => n17400, ZN => n17570);
   U13014 : NOR2_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_0_port, A2
                           => n13876, ZN => n17571);
   U13015 : NAND2_X1 port map( A1 => n17663, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_0_port, ZN => n17574);
   U13016 : NOR2_X1 port map( A1 => pipeline_EXE_controls_in_EXEcute_0_port, A2
                           => n13848, ZN => n17577);
   U13017 : NOR2_X1 port map( A1 => n17667, A2 => n17397, ZN => n17552);
   U13018 : AOI221_X1 port map( B1 => n17340, B2 => 
                           pipeline_Reg1_Addr_to_exe_3_port, C1 => 
                           pipeline_regDst_to_mem_4_port, C2 => n17399, A => 
                           n16811, ZN => n16806);
   U13019 : NOR4_X1 port map( A1 => n17559, A2 => n17560, A3 => n17561, A4 => 
                           n17562, ZN => n17557);
   U13020 : OAI21_X1 port map( B1 => n17385, B2 => 
                           pipeline_Reg1_Addr_to_exe_3_port, A => n17563, ZN =>
                           n17562);
   U13021 : NAND2_X1 port map( A1 => n17386, A2 => 
                           pipeline_Reg1_Addr_to_exe_4_port, ZN => n17563);
   U13022 : OAI21_X1 port map( B1 => n17314, B2 => 
                           pipeline_Reg1_Addr_to_exe_0_port, A => n17564, ZN =>
                           n17561);
   U13023 : NAND2_X1 port map( A1 => n17385, A2 => 
                           pipeline_Reg1_Addr_to_exe_3_port, ZN => n17564);
   U13024 : OAI21_X1 port map( B1 => pipeline_Reg1_Addr_to_exe_1_port, B2 => 
                           n17304, A => n17565, ZN => n17560);
   U13025 : NAND2_X1 port map( A1 => n17314, A2 => 
                           pipeline_Reg1_Addr_to_exe_0_port, ZN => n17565);
   U13026 : OAI211_X1 port map( C1 => n17386, C2 => 
                           pipeline_Reg1_Addr_to_exe_4_port, A => n17566, B => 
                           n17567, ZN => n17559);
   U13027 : NAND2_X1 port map( A1 => n17304, A2 => 
                           pipeline_Reg1_Addr_to_exe_1_port, ZN => n17566);
   U13028 : NAND2_X1 port map( A1 => n17333, A2 => 
                           pipeline_data_to_RF_from_WB_30_port, ZN => n17639);
   U13029 : NAND2_X1 port map( A1 => n17106, A2 => n17640, ZN => n17637);
   U13030 : NOR2_X1 port map( A1 => n15834, A2 => n14127, ZN => n17675);
   U13031 : NOR2_X1 port map( A1 => n16529, A2 => n16528, ZN => n17345);
   U13032 : NOR2_X1 port map( A1 => n16529, A2 => n16528, ZN => n17337);
   U13033 : NOR2_X1 port map( A1 => n16530, A2 => n16531, ZN => n17339);
   U13034 : NOR2_X1 port map( A1 => n16533, A2 => n16532, ZN => n17335);
   U13035 : NOR2_X1 port map( A1 => n16527, A2 => n16539, ZN => n17342);
   U13036 : NOR2_X1 port map( A1 => n16529, A2 => n16528, ZN => n17336);
   U13037 : NOR2_X1 port map( A1 => n16530, A2 => n16531, ZN => n17338);
   U13038 : NOR2_X1 port map( A1 => n16533, A2 => n16532, ZN => n17334);
   U13039 : NOR2_X1 port map( A1 => n16527, A2 => n16539, ZN => n17341);
   U13040 : OAI221_X1 port map( B1 => pipeline_RegDst_to_WB_2_port, B2 => 
                           n17383, C1 => n17326, C2 => 
                           pipeline_stageD_offset_jump_sign_ext_23_port, A => 
                           n16565, ZN => n16563);
   U13041 : AOI221_X1 port map( B1 => pipeline_regDst_to_mem_3_port, B2 => 
                           n17384, C1 => n17340, C2 => 
                           pipeline_stageD_offset_jump_sign_ext_24_port, A => 
                           n16573, ZN => n16572);
   U13042 : NOR2_X1 port map( A1 => n14879, A2 => n14860, ZN => n14245);
   U13043 : NOR2_X1 port map( A1 => n14879, A2 => n14864, ZN => n14239);
   U13044 : NOR2_X1 port map( A1 => n14860, A2 => n14873, ZN => n14227);
   U13045 : NOR2_X1 port map( A1 => n14863, A2 => n14867, ZN => n14224);
   U13046 : NOR3_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_add_alu_sCout_0_port, A2 => 
                           pipeline_EXE_controls_in_EXEcute_2_port, A3 => 
                           n15586, ZN => n14965);
   U13047 : NOR2_X1 port map( A1 => n14878, A2 => n14860, ZN => n14246);
   U13048 : NOR2_X1 port map( A1 => n15348, A2 => 
                           pipeline_stageE_input1_to_ALU_18_port, ZN => n16631)
                           ;
   U13049 : NOR2_X1 port map( A1 => n14865, A2 => n14866, ZN => n14225);
   U13050 : NOR2_X1 port map( A1 => n14864, A2 => n14866, ZN => n14222);
   U13051 : NOR2_X1 port map( A1 => n14865, A2 => n14872, ZN => n14236);
   U13052 : NOR2_X1 port map( A1 => n14864, A2 => n14872, ZN => n14234);
   U13053 : NOR2_X1 port map( A1 => n14860, A2 => n14872, ZN => n14228);
   U13054 : NOR2_X1 port map( A1 => n14865, A2 => n14862, ZN => n14244);
   U13055 : NOR3_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_add_alu_sCout_0_port, A2 => 
                           n17405, A3 => n15586, ZN => n14966);
   U13056 : NOR2_X1 port map( A1 => n16609, A2 => 
                           pipeline_stageE_input1_to_ALU_29_port, ZN => n15164)
                           ;
   U13057 : NAND2_X1 port map( A1 => pipeline_stageE_EXE_ALU_alu_shift_N202, A2
                           => n14961, ZN => n17429);
   U13058 : NAND4_X1 port map( A1 => n17609, A2 => n17610, A3 => n17611, A4 => 
                           n15163, ZN => n17541);
   U13059 : NAND2_X1 port map( A1 => n17636, A2 => n17402, ZN => n3989);
   U13060 : NOR2_X1 port map( A1 => n17537, A2 => n17538, ZN => n17536);
   U13061 : NAND2_X1 port map( A1 => n17535, A2 => n17536, ZN => n17534);
   U13062 : NOR3_X1 port map( A1 => n15014, A2 => n15013, A3 => n17534, ZN => 
                           n17533);
   U13063 : AOI21_X1 port map( B1 => n17539, B2 => n17615, A => n17616, ZN => 
                           n17613);
   U13064 : XNOR2_X1 port map( A => n17539, B => n15191, ZN => n15011);
   U13065 : OAI21_X1 port map( B1 => n17539, B2 => n15146, A => n15145, ZN => 
                           n15159);
   U13066 : NAND2_X1 port map( A1 => n17541, A2 => n15166, ZN => n17544);
   U13067 : NAND2_X1 port map( A1 => n17541, A2 => n17540, ZN => n17543);
   U13068 : NAND2_X1 port map( A1 => n17543, A2 => n15147, ZN => n17542);
   U13069 : XNOR2_X1 port map( A => n17544, B => n17612, ZN => n15010);
   U13070 : NAND3_X1 port map( A1 => n15010, A2 => n15009, A3 => n17546, ZN => 
                           n17545);
   U13071 : NAND2_X1 port map( A1 => n17547, A2 => n17551, ZN => n17619);
   U13072 : NOR2_X1 port map( A1 => n17545, A2 => n17550, ZN => n17620);
   U13073 : OAI211_X1 port map( C1 => n17542, C2 => n15161, A => n15142, B => 
                           n13939, ZN => n16598);
   U13074 : OAI22_X1 port map( A1 => n17314, A2 => 
                           pipeline_Reg2_Addr_to_exe_0_port, B1 => n17385, B2 
                           => pipeline_Reg2_Addr_to_exe_3_port, ZN => n16783);
   U13075 : NOR3_X1 port map( A1 => n17548, A2 => n17549, A3 => n16783, ZN => 
                           n16782);
   U13076 : OAI221_X1 port map( B1 => pipeline_RegDst_to_WB_2_port, B2 => 
                           n17403, C1 => n17326, C2 => 
                           pipeline_Reg2_Addr_to_exe_2_port, A => n16782, ZN =>
                           n16780);
   U13077 : NAND2_X1 port map( A1 => n17411, A2 => n17551, ZN => n17550);
   U13078 : AOI21_X1 port map( B1 => n17619, B2 => n17618, A => n17620, ZN => 
                           n15000);
   U13079 : AOI21_X1 port map( B1 => n16584, B2 => n16805, A => n13940, ZN => 
                           n16585);
   U13080 : AOI21_X1 port map( B1 => n15123, B2 => 
                           pipeline_data_to_RF_from_WB_1_port, A => n17552, ZN 
                           => n16699);
   U13081 : OAI22_X1 port map( A1 => n17393, A2 => 
                           pipeline_Reg2_Addr_to_exe_4_port, B1 => n17340, B2 
                           => pipeline_Reg2_Addr_to_exe_3_port, ZN => n17555);
   U13082 : AOI22_X1 port map( A1 => n17393, A2 => 
                           pipeline_Reg2_Addr_to_exe_4_port, B1 => n17340, B2 
                           => pipeline_Reg2_Addr_to_exe_3_port, ZN => n17554);
   U13083 : NAND2_X1 port map( A1 => n17553, A2 => n17554, ZN => n16786);
   U13084 : NOR4_X1 port map( A1 => n16561, A2 => n16780, A3 => n16779, A4 => 
                           n16778, ZN => n17668);
   U13085 : NOR2_X1 port map( A1 => n17667, A2 => n17398, ZN => n17556);
   U13086 : AOI21_X1 port map( B1 => n17669, B2 => 
                           pipeline_data_to_RF_from_WB_2_port, A => n17556, ZN 
                           => n16704);
   U13087 : NAND3_X1 port map( A1 => n17643, A2 => n17557, A3 => n17558, ZN => 
                           n16617);
   U13088 : XOR2_X1 port map( A => n17401, B => pipeline_RegDst_to_WB_2_port, Z
                           => n17567);
   U13089 : NAND2_X1 port map( A1 => n17642, A2 => n16696, ZN => n17568);
   U13090 : NAND2_X1 port map( A1 => n16696, A2 => n17571, ZN => n17569);
   U13091 : OAI21_X1 port map( B1 => n17666, B2 => n17123, A => n17327, ZN => 
                           n17641);
   U13092 : OAI21_X1 port map( B1 => n17105, B2 => n17396, A => n17574, ZN => 
                           n17573);
   U13093 : AOI21_X1 port map( B1 => n17073, B2 => 
                           pipeline_stageE_EXE_ALU_add_alu_sCout_0_port, A => 
                           n17576, ZN => n16691);
   U13094 : OAI22_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_1_port, A2 
                           => n17381, B1 => n17741, B2 => 
                           pipeline_stageE_EXE_ALU_add_alu_sCout_0_port, ZN => 
                           n16693);
   U13095 : NAND2_X1 port map( A1 => n15049, A2 => n15048, ZN => n17578);
   U13096 : NAND2_X1 port map( A1 => n15050, A2 => n17578, ZN => n16690);
   U13097 : OAI21_X1 port map( B1 => n15055, B2 => n16690, A => n15053, ZN => 
                           n16688);
   U13098 : OAI21_X1 port map( B1 => n15055, B2 => n16690, A => n15053, ZN => 
                           n17579);
   U13099 : NAND2_X1 port map( A1 => n15566, A2 => n15569, ZN => n16682);
   U13100 : NAND2_X1 port map( A1 => n16682, A2 => n15568, ZN => n15541);
   U13101 : NAND3_X1 port map( A1 => n17582, A2 => n15527, A3 => n17583, ZN => 
                           n17580);
   U13102 : OAI21_X1 port map( B1 => n15541, B2 => n15542, A => n17584, ZN => 
                           n17582);
   U13103 : NAND2_X1 port map( A1 => n17580, A2 => n17581, ZN => n15508);
   U13104 : NAND2_X1 port map( A1 => n15508, A2 => n15509, ZN => n15478);
   U13105 : NAND3_X1 port map( A1 => n17585, A2 => n15463, A3 => n17586, ZN => 
                           n16664);
   U13106 : NAND3_X1 port map( A1 => n15494, A2 => n15495, A3 => n17587, ZN => 
                           n17585);
   U13107 : NAND2_X1 port map( A1 => n16664, A2 => 
                           pipeline_stageE_input1_to_ALU_11_port, ZN => n17588)
                           ;
   U13108 : NAND2_X1 port map( A1 => n16664, A2 => n15459, ZN => n17589);
   U13109 : NAND3_X1 port map( A1 => n15367, A2 => n15383, A3 => n16630, ZN => 
                           n17601);
   U13110 : NAND2_X1 port map( A1 => n15368, A2 => n17600, ZN => n17593);
   U13111 : OAI221_X1 port map( B1 => n15248, B2 => n17117, C1 => n15248, C2 =>
                           n16613, A => n15250, ZN => n15235);
   U13112 : XOR2_X1 port map( A => n17078, B => n15204, Z => n17607);
   U13113 : XNOR2_X1 port map( A => n15205, B => n17607, ZN => n15014);
   U13114 : NAND2_X1 port map( A1 => n15205, A2 => 
                           pipeline_stageE_input1_to_ALU_27_port, ZN => n17609)
                           ;
   U13115 : NAND2_X1 port map( A1 => n15205, A2 => n15204, ZN => n17610);
   U13116 : XNOR2_X1 port map( A => n17613, B => n17614, ZN => n15007);
   U13117 : OAI211_X1 port map( C1 => n15046, C2 => n14949, A => n17429, B => 
                           n17629, ZN => n17628);
   U13118 : AOI21_X1 port map( B1 => pipeline_stageE_EXE_ALU_alu_shift_N234, B2
                           => n17681, A => n17628, ZN => n17627);
   U13119 : NAND2_X1 port map( A1 => pipeline_stageE_EXE_ALU_alu_shift_N39, A2 
                           => n17149, ZN => n17626);
   U13120 : NAND2_X1 port map( A1 => n17624, A2 => n17635, ZN => n17623);
   U13121 : NAND2_X1 port map( A1 => n17630, A2 => n14995, ZN => n17629);
   U13122 : NAND2_X1 port map( A1 => pipeline_stageE_EXE_ALU_alu_shift_N7, A2 
                           => n14965, ZN => n17625);
   U13123 : NAND2_X1 port map( A1 => pipeline_stageE_EXE_ALU_alu_shift_N137, A2
                           => n17680, ZN => n17624);
   U13124 : NAND2_X1 port map( A1 => pipeline_stageD_target_Jump_temp_30_port, 
                           A2 => n17675, ZN => n17636);
   U13125 : OAI221_X1 port map( B1 => 
                           pipeline_stageD_offset_to_jump_temp_7_port, B2 => 
                           pipeline_stageD_offset_to_jump_temp_2_port, C1 => 
                           pipeline_stageD_offset_to_jump_temp_7_port, C2 => 
                           n17406, A => pipeline_cu_pipeline_N89, ZN => n14072)
                           ;
   U13126 : NOR4_X1 port map( A1 => pipeline_stageD_offset_to_jump_temp_3_port,
                           A2 => pipeline_stageD_offset_to_jump_temp_4_port, A3
                           => pipeline_stageD_offset_to_jump_temp_2_port, A4 =>
                           n17350, ZN => n13990);
   U13127 : AOI22_X1 port map( A1 => n17671, A2 => 
                           pipeline_stageD_offset_to_jump_temp_2_port, B1 => 
                           n17107, B2 => InstrFetched_2_port, ZN => n15623);
   U13128 : NAND4_X1 port map( A1 => pipeline_stageD_offset_to_jump_temp_3_port
                           , A2 => pipeline_stageD_offset_to_jump_temp_5_port, 
                           A3 => pipeline_stageD_offset_to_jump_temp_2_port, A4
                           => n17406, ZN => n14180);
   U13129 : NOR3_X1 port map( A1 => pipeline_stageD_offset_to_jump_temp_2_port,
                           A2 => n17410, A3 => n17350, ZN => n14179);
   U13130 : AOI22_X1 port map( A1 => n17671, A2 => 
                           pipeline_nextPC_IFID_DEC_0_port, B1 => n17673, B2 =>
                           pipeline_stageF_PC_plus4_N7, ZN => n15773);
   U13131 : AOI22_X1 port map( A1 => n17663, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_29_port, B1 => n16620, 
                           B2 => n13956, ZN => n16770);
   U13132 : AOI22_X1 port map( A1 => n17663, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_28_port, B1 => n16620, 
                           B2 => n13962, ZN => n16766);
   U13133 : AOI22_X1 port map( A1 => n17663, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_23_port, B1 => n16620, 
                           B2 => n13952, ZN => n16753);
   U13134 : AOI22_X1 port map( A1 => n17663, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_19_port, B1 => n16620, 
                           B2 => n13948, ZN => n16637);
   U13135 : AOI22_X1 port map( A1 => n17663, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_15_port, B1 => n16620, 
                           B2 => n13959, ZN => n16733);
   U13136 : AOI22_X1 port map( A1 => n17663, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_18_port, B1 => n16620, 
                           B2 => n13947, ZN => n16734);
   U13137 : AOI22_X1 port map( A1 => n17663, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_16_port, B1 => n16620, 
                           B2 => n13804, ZN => n16641);
   U13138 : AOI22_X1 port map( A1 => n17663, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_9_port, B1 => n16620, 
                           B2 => n13820, ZN => n16671);
   U13139 : AOI22_X1 port map( A1 => n17663, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_8_port, B1 => n16620, 
                           B2 => n13964, ZN => n16720);
   U13140 : AOI22_X1 port map( A1 => n17663, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_1_port, B1 => n16620, 
                           B2 => n13847, ZN => n16701);
   U13141 : XNOR2_X1 port map( A => 
                           pipeline_stageE_EXE_ALU_add_alu_sCout_0_port, B => 
                           n15133, ZN => n15137);
   U13142 : XNOR2_X1 port map( A => n15493, B => n15494, ZN => n15035);
   U13143 : OAI221_X1 port map( B1 => n15477, B2 => n15478, C1 => n15477, C2 =>
                           n15479, A => n15480, ZN => n15476);
   U13144 : AOI22_X1 port map( A1 => n17665, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_29_port, B1 => n17123, 
                           B2 => pipeline_data_to_RF_from_WB_29_port, ZN => 
                           n16773);
   U13145 : AOI22_X1 port map( A1 => n17666, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_25_port, B1 => n17123, 
                           B2 => pipeline_data_to_RF_from_WB_25_port, ZN => 
                           n16757);
   U13146 : AOI22_X1 port map( A1 => n17666, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_23_port, B1 => n17123, 
                           B2 => pipeline_data_to_RF_from_WB_23_port, ZN => 
                           n16752);
   U13147 : AOI22_X1 port map( A1 => n17666, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_16_port, B1 => n17123, 
                           B2 => pipeline_data_to_RF_from_WB_16_port, ZN => 
                           n16640);
   U13148 : AOI22_X1 port map( A1 => n17665, A2 => 
                           pipeline_Alu_Out_Addr_to_mem_12_port, B1 => n17123, 
                           B2 => pipeline_data_to_RF_from_WB_12_port, ZN => 
                           n16663);
   U13149 : NOR2_X1 port map( A1 => n17340, A2 => n14129, ZN => 
                           pipeline_MEMWB_Stage_N46);
   U13150 : OAI22_X1 port map( A1 => n17304, A2 => 
                           pipeline_stageD_offset_jump_sign_ext_22_port, B1 => 
                           n17386, B2 => 
                           pipeline_stageD_offset_jump_sign_ext_31_port, ZN => 
                           n16568);
   U13151 : AOI22_X1 port map( A1 => n17304, A2 => 
                           pipeline_Reg2_Addr_to_exe_1_port, B1 => 
                           pipeline_Reg2_Addr_to_exe_4_port, B2 => n17386, ZN 
                           => n16784);
   U13152 : NAND3_X1 port map( A1 => n15368, A2 => n15367, A3 => n15383, ZN => 
                           n17648);
   U13153 : AOI22_X1 port map( A1 => pipeline_data_to_RF_from_WB_0_port, A2 => 
                           n17123, B1 => pipeline_Alu_Out_Addr_to_mem_0_port, 
                           B2 => n17665, ZN => n16696);
   U13154 : OAI21_X1 port map( B1 => n15596, B2 => 
                           pipeline_stageE_EXE_ALU_alu_shift_N202, A => n15050,
                           ZN => n15597);
   U13155 : NOR2_X1 port map( A1 => n16631, A2 => n17648, ZN => n17649);
   U13156 : NAND2_X1 port map( A1 => n15049, A2 => n15050, ZN => n15047);
   U13157 : NAND2_X1 port map( A1 => n16806, A2 => n16807, ZN => n16796);
   U13158 : NAND2_X1 port map( A1 => n15049, A2 => n15595, ZN => n15056);
   U13159 : NOR4_X1 port map( A1 => n16778, A2 => n16561, A3 => n16779, A4 => 
                           n16780, ZN => n15123);
   U13160 : XNOR2_X1 port map( A => n15554, B => n15541, ZN => n15042);
   U13161 : AOI21_X1 port map( B1 => n15540, B2 => n15541, A => n15542, ZN => 
                           n15526);
   U13162 : NOR2_X1 port map( A1 => n16554, A2 => n16555, ZN => n14103);
   U13163 : OAI221_X1 port map( B1 => pipeline_regDst_to_mem_4_port, B2 => 
                           n17328, C1 => n17393, C2 => 
                           pipeline_stageD_offset_jump_sign_ext_31_port, A => 
                           n16574, ZN => n16573);
   U13164 : OAI22_X1 port map( A1 => n17340, A2 => 
                           pipeline_Reg1_Addr_to_exe_3_port, B1 => n17399, B2 
                           => pipeline_regDst_to_mem_4_port, ZN => n16811);
   U13165 : OAI22_X1 port map( A1 => pipeline_stageE_EXE_ALU_alu_shift_N202, A2
                           => pipeline_stageE_EXE_ALU_alu_shift_C48_SH_0_port, 
                           B1 => n17742, B2 => n17119, ZN => n15046);
   U13166 : AOI22_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_add_alu_sCout_0_port, A2 => 
                           pipeline_stageE_input2_to_ALU_0_port, B1 => n17742, 
                           B2 => n17381, ZN => n15596);
   U13167 : AOI21_X1 port map( B1 => n15416, B2 => n16652, A => n15413, ZN => 
                           n16650);
   U13168 : OAI211_X1 port map( C1 => net175543, C2 => n13990, A => 
                           pipeline_stageD_offset_to_jump_temp_1_port, B => 
                           pipeline_cu_pipeline_N89, ZN => n14071);
   U13169 : AOI22_X1 port map( A1 => n17671, A2 => net175543, B1 => n15601, B2 
                           => InstrFetched_0_port, ZN => n15621);
   U13170 : NOR2_X1 port map( A1 => net175543, A2 => n17406, ZN => n14051);
   U13171 : NOR2_X1 port map( A1 => pipeline_stageD_offset_to_jump_temp_1_port,
                           A2 => net175543, ZN => n14032);
   U13172 : XNOR2_X1 port map( A => n15047, B => n15048, ZN => n14970);
   U13173 : NOR3_X1 port map( A1 => 
                           pipeline_stageE_EXE_ALU_alu_shift_C48_SH_1_port, A2 
                           => pipeline_stageE_input1_to_ALU_1_port, A3 => 
                           n17678, ZN => n14974);
   U13174 : AOI211_X1 port map( C1 => n14993, C2 => n15007, A => n15126, B => 
                           n15127, ZN => n15125);
   U13175 : XNOR2_X1 port map( A => n15217, B => n15218, ZN => n15015);
   U13176 : XNOR2_X1 port map( A => n15234, B => n15235, ZN => n15233);
   U13177 : NAND2_X1 port map( A1 => n15445, A2 => n15446, ZN => n16657);
   U13178 : NOR2_X1 port map( A1 => n16650, A2 => n15398, ZN => n16646);

end SYN_struct;
